module mod0 #(parameter KRATOS_INSTANCE_ID = 32'h0)
(
    input I
);

endmodule   // mod
