module Main (
    input [4:0] I [4:0],
    output [4:0] O [4:0]
);
wire [24:0] x;
assign x = {I[4][4],I[4][3],I[4][2],I[4][1],I[4][0],I[3][4],I[3][3],I[3][2],I[3][1],I[3][0],I[2][4],I[2][3],I[2][2],I[2][1],I[2][0],I[1][4],I[1][3],I[1][2],I[1][1],I[1][0],I[0][4],I[0][3],I[0][2],I[0][1],I[0][0]};
assign O[4] = {x[24],x[23],x[22],x[21],x[20]};
assign O[3] = {x[19],x[18],x[17],x[16],x[15]};
assign O[2] = {x[14],x[13],x[12],x[11],x[10]};
assign O[1] = {x[9],x[8],x[7],x[6],x[5]};
assign O[0] = {x[4],x[3],x[2],x[1],x[0]};
endmodule

