module return_magma_tuple (input [1:0] I_0, output  O_0, output  O_1);
assign O_0 = I_0[0];
assign O_1 = I_0[1];
endmodule

