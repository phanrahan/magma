module test_reduce_xor (
    input [4:0] I,
    output O
);
assign O = ^ I;
endmodule

