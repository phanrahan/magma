module Test (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

