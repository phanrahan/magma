module no_outputs(	// <stdin>:1:1
  input I);

endmodule

