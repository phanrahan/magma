module Main (
    output [3:0][4:0][2:0] a0,
    output [3:0][4:0][2:0] a1,
    input [3:0][4:0][1:0] b,
    input [2:0][1:0] c
);
assign a0 = {{{1'b0,1'b0,1'b0},{1'b0,1'b0,1'b0},{1'b0,1'b0,1'b0},{1'b0,1'b0,1'b0},{1'b0,1'b0,1'b0}},{{1'b0,1'b0,1'b0},{1'b0,1'b0},b[1][4],b[1][3]},{b[1][2],b[1][1],b[1][0],b[0][4]},{b[0][3],b[0][2],b[0][1],b[0][0]}};
assign a1 = {{{1'b0,1'b0,1'b0},{1'b0,1'b0,1'b0},{1'b0,1'b0,1'b0},{1'b0,1'b0,1'b0},{1'b0,1'b0,1'b0}},{{1'b0,1'b0,1'b0},{1'b0,1'b0,1'b0},{c[1][2],1'b0,1'b0},{1'b0,c[1][1],1'b0},{1'b0,1'b0,c[1][0]}},{{1'b0,1'b0,1'b0},{1'b0,1'b0,1'b0},{1'b0,1'b0,1'b0},{1'b0,1'b0,c[0][2]},{1'b0,1'b0,1'b0}},{{c[0][1],1'b0,1'b0},{1'b0,c[0][0],1'b0},{1'b0,1'b0,1'b0},{1'b0,1'b0,1'b0},{1'b0,1'b0,1'b0}}};
endmodule

