module Main (
    input I,
    output O0,
    output O1
);
wire x;
assign x = I;
assign O0 = x;
assign O1 = x;
endmodule

