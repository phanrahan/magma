module mod1 #(parameter KRATOS_INSTANCE_ID = 'hEF)
(
    input I
);

endmodule   // mod
