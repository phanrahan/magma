module coreir_term #(
    parameter width = 1
) (
    input [width-1:0] in
);

endmodule

module MonitorWrapper (
    input [7:0] arr [63:0]
);
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_1;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_2;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_3;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_4;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_5;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_6;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_7;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_8;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_9;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_10;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_11;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_12;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_13;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_14;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_15;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_16;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_17;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_18;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_19;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_20;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_21;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_22;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_23;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_24;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_25;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_26;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_27;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_28;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_29;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_30;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_31;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_32;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_33;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_34;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_35;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_36;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_37;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_38;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_39;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_40;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_41;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_42;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_43;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_44;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_45;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_46;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_47;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_48;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_49;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_50;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_51;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_52;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_53;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_54;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_55;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_56;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_57;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_58;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_59;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_60;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_61;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_62;
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_63;
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0 = arr[63];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_1 = arr[62];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_2 = arr[61];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_3 = arr[60];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_4 = arr[59];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_5 = arr[58];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_6 = arr[57];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_7 = arr[56];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_8 = arr[55];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_9 = arr[54];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_10 = arr[53];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_11 = arr[52];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_12 = arr[51];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_13 = arr[50];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_14 = arr[49];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_15 = arr[48];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_16 = arr[47];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_17 = arr[46];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_18 = arr[45];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_19 = arr[44];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_20 = arr[43];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_21 = arr[42];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_22 = arr[41];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_23 = arr[40];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_24 = arr[39];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_25 = arr[38];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_26 = arr[37];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_27 = arr[36];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_28 = arr[35];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_29 = arr[34];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_30 = arr[33];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_31 = arr[32];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_32 = arr[31];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_33 = arr[30];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_34 = arr[29];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_35 = arr[28];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_36 = arr[27];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_37 = arr[26];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_38 = arr[25];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_39 = arr[24];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_40 = arr[23];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_41 = arr[22];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_42 = arr[21];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_43 = arr[20];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_44 = arr[19];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_45 = arr[18];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_46 = arr[17];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_47 = arr[16];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_48 = arr[15];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_49 = arr[14];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_50 = arr[13];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_51 = arr[12];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_52 = arr[11];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_53 = arr[10];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_54 = arr[9];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_55 = arr[8];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_56 = arr[7];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_57 = arr[6];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_58 = arr[5];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_59 = arr[4];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_60 = arr[3];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_61 = arr[2];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_62 = arr[1];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_63 = arr[0];

monitor #(.WIDTH(8), .DEPTH(64)) monitor_inst(.arr('{MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_1, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_2, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_3, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_4, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_5, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_6, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_7, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_8, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_9, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_10, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_11, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_12, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_13, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_14, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_15, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_16, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_17, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_18, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_19, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_20, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_21, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_22, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_23, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_24, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_25, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_26, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_27, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_28, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_29, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_30, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_31, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_32, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_33, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_34, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_35, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_36, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_37, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_38, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_39, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_40, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_41, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_42, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_43, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_44, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_45, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_46, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_47, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_48, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_49, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_50, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_51, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_52, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_53, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_54, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_55, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_56, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_57, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_58, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_59, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_60, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_61, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_62, MonitorWrapper_inline_verilog_inst_0___magma_inline_value_63}));
                    
endmodule

