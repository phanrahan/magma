module simple_inline_verilog2(
  input  I,
  output O
);


  	// This is 'a' "comment".
  assign O = I;
endmodule

