module top(a, b);
    input a;
    output b;
    assign a = b;
endmodule
