module file(
  input                                                        CLK, ASYNCRESET,
  input  [7:0]                                                 file_read_0_addr,
  input  [7:0]                                                 file_read_1_addr,
  input  struct packed {logic [31:0] data; logic [7:0] addr; } write_0,
  input                                                        write_0_en,
  output [31:0]                                                file_read_0_data,
  output [31:0]                                                file_read_1_data);

  reg [31:0] Register_inst0;
  reg [31:0] Register_inst1;
  reg [31:0] Register_inst2;
  reg [31:0] Register_inst3;
  reg [31:0] Register_inst4;
  reg [31:0] Register_inst5;
  reg [31:0] Register_inst6;
  reg [31:0] Register_inst7;
  reg [31:0] Register_inst8;
  reg [31:0] Register_inst9;
  reg [31:0] Register_inst10;
  reg [31:0] Register_inst11;
  reg [31:0] Register_inst12;
  reg [31:0] Register_inst13;
  reg [31:0] Register_inst14;
  reg [31:0] Register_inst15;
  reg [31:0] Register_inst16;
  reg [31:0] Register_inst17;
  reg [31:0] Register_inst18;
  reg [31:0] Register_inst19;
  reg [31:0] Register_inst20;
  reg [31:0] Register_inst21;
  reg [31:0] Register_inst22;
  reg [31:0] Register_inst23;
  reg [31:0] Register_inst24;
  reg [31:0] Register_inst25;
  reg [31:0] Register_inst26;
  reg [31:0] Register_inst27;
  reg [31:0] Register_inst28;
  reg [31:0] Register_inst29;
  reg [31:0] Register_inst30;
  reg [31:0] Register_inst31;
  reg [31:0] Register_inst32;
  reg [31:0] Register_inst33;
  reg [31:0] Register_inst34;
  reg [31:0] Register_inst35;
  reg [31:0] Register_inst36;
  reg [31:0] Register_inst37;
  reg [31:0] Register_inst38;
  reg [31:0] Register_inst39;
  reg [31:0] Register_inst40;
  reg [31:0] Register_inst41;
  reg [31:0] Register_inst42;
  reg [31:0] Register_inst43;
  reg [31:0] Register_inst44;
  reg [31:0] Register_inst45;
  reg [31:0] Register_inst46;
  reg [31:0] Register_inst47;
  reg [31:0] Register_inst48;
  reg [31:0] Register_inst49;
  reg [31:0] Register_inst50;
  reg [31:0] Register_inst51;
  reg [31:0] Register_inst52;
  reg [31:0] Register_inst53;
  reg [31:0] Register_inst54;
  reg [31:0] Register_inst55;
  reg [31:0] Register_inst56;
  reg [31:0] Register_inst57;
  reg [31:0] Register_inst58;
  reg [31:0] Register_inst59;
  reg [31:0] Register_inst60;
  reg [31:0] Register_inst61;
  reg [31:0] Register_inst62;
  reg [31:0] Register_inst63;
  reg [31:0] Register_inst64;
  reg [31:0] Register_inst65;
  reg [31:0] Register_inst66;
  reg [31:0] Register_inst67;
  reg [31:0] Register_inst68;
  reg [31:0] Register_inst69;
  reg [31:0] Register_inst70;
  reg [31:0] Register_inst71;
  reg [31:0] Register_inst72;
  reg [31:0] Register_inst73;
  reg [31:0] Register_inst74;
  reg [31:0] Register_inst75;
  reg [31:0] Register_inst76;
  reg [31:0] Register_inst77;
  reg [31:0] Register_inst78;
  reg [31:0] Register_inst79;
  reg [31:0] Register_inst80;
  reg [31:0] Register_inst81;
  reg [31:0] Register_inst82;
  reg [31:0] Register_inst83;
  reg [31:0] Register_inst84;
  reg [31:0] Register_inst85;
  reg [31:0] Register_inst86;
  reg [31:0] Register_inst87;
  reg [31:0] Register_inst88;
  reg [31:0] Register_inst89;
  reg [31:0] Register_inst90;
  reg [31:0] Register_inst91;
  reg [31:0] Register_inst92;
  reg [31:0] Register_inst93;
  reg [31:0] Register_inst94;
  reg [31:0] Register_inst95;
  reg [31:0] Register_inst96;
  reg [31:0] Register_inst97;
  reg [31:0] Register_inst98;
  reg [31:0] Register_inst99;
  reg [31:0] Register_inst100;
  reg [31:0] Register_inst101;
  reg [31:0] Register_inst102;
  reg [31:0] Register_inst103;
  reg [31:0] Register_inst104;
  reg [31:0] Register_inst105;
  reg [31:0] Register_inst106;
  reg [31:0] Register_inst107;
  reg [31:0] Register_inst108;
  reg [31:0] Register_inst109;
  reg [31:0] Register_inst110;
  reg [31:0] Register_inst111;
  reg [31:0] Register_inst112;
  reg [31:0] Register_inst113;
  reg [31:0] Register_inst114;
  reg [31:0] Register_inst115;
  reg [31:0] Register_inst116;
  reg [31:0] Register_inst117;
  reg [31:0] Register_inst118;
  reg [31:0] Register_inst119;
  reg [31:0] Register_inst120;
  reg [31:0] Register_inst121;
  reg [31:0] Register_inst122;
  reg [31:0] Register_inst123;
  reg [31:0] Register_inst124;
  reg [31:0] Register_inst125;
  reg [31:0] Register_inst126;
  reg [31:0] Register_inst127;
  reg [31:0] Register_inst128;
  reg [31:0] Register_inst129;
  reg [31:0] Register_inst130;
  reg [31:0] Register_inst131;
  reg [31:0] Register_inst132;
  reg [31:0] Register_inst133;
  reg [31:0] Register_inst134;
  reg [31:0] Register_inst135;
  reg [31:0] Register_inst136;
  reg [31:0] Register_inst137;
  reg [31:0] Register_inst138;
  reg [31:0] Register_inst139;
  reg [31:0] Register_inst140;
  reg [31:0] Register_inst141;
  reg [31:0] Register_inst142;
  reg [31:0] Register_inst143;
  reg [31:0] Register_inst144;
  reg [31:0] Register_inst145;
  reg [31:0] Register_inst146;
  reg [31:0] Register_inst147;
  reg [31:0] Register_inst148;
  reg [31:0] Register_inst149;
  reg [31:0] Register_inst150;
  reg [31:0] Register_inst151;
  reg [31:0] Register_inst152;
  reg [31:0] Register_inst153;
  reg [31:0] Register_inst154;
  reg [31:0] Register_inst155;
  reg [31:0] Register_inst156;
  reg [31:0] Register_inst157;
  reg [31:0] Register_inst158;
  reg [31:0] Register_inst159;
  reg [31:0] Register_inst160;
  reg [31:0] Register_inst161;
  reg [31:0] Register_inst162;
  reg [31:0] Register_inst163;
  reg [31:0] Register_inst164;
  reg [31:0] Register_inst165;
  reg [31:0] Register_inst166;
  reg [31:0] Register_inst167;
  reg [31:0] Register_inst168;
  reg [31:0] Register_inst169;
  reg [31:0] Register_inst170;
  reg [31:0] Register_inst171;
  reg [31:0] Register_inst172;
  reg [31:0] Register_inst173;
  reg [31:0] Register_inst174;
  reg [31:0] Register_inst175;
  reg [31:0] Register_inst176;
  reg [31:0] Register_inst177;
  reg [31:0] Register_inst178;
  reg [31:0] Register_inst179;
  reg [31:0] Register_inst180;
  reg [31:0] Register_inst181;
  reg [31:0] Register_inst182;
  reg [31:0] Register_inst183;
  reg [31:0] Register_inst184;
  reg [31:0] Register_inst185;
  reg [31:0] Register_inst186;
  reg [31:0] Register_inst187;
  reg [31:0] Register_inst188;
  reg [31:0] Register_inst189;
  reg [31:0] Register_inst190;
  reg [31:0] Register_inst191;
  reg [31:0] Register_inst192;
  reg [31:0] Register_inst193;
  reg [31:0] Register_inst194;
  reg [31:0] Register_inst195;
  reg [31:0] Register_inst196;
  reg [31:0] Register_inst197;
  reg [31:0] Register_inst198;
  reg [31:0] Register_inst199;
  reg [31:0] Register_inst200;
  reg [31:0] Register_inst201;
  reg [31:0] Register_inst202;
  reg [31:0] Register_inst203;
  reg [31:0] Register_inst204;
  reg [31:0] Register_inst205;
  reg [31:0] Register_inst206;
  reg [31:0] Register_inst207;
  reg [31:0] Register_inst208;
  reg [31:0] Register_inst209;
  reg [31:0] Register_inst210;
  reg [31:0] Register_inst211;
  reg [31:0] Register_inst212;
  reg [31:0] Register_inst213;
  reg [31:0] Register_inst214;
  reg [31:0] Register_inst215;
  reg [31:0] Register_inst216;
  reg [31:0] Register_inst217;
  reg [31:0] Register_inst218;
  reg [31:0] Register_inst219;
  reg [31:0] Register_inst220;
  reg [31:0] Register_inst221;
  reg [31:0] Register_inst222;
  reg [31:0] Register_inst223;
  reg [31:0] Register_inst224;
  reg [31:0] Register_inst225;
  reg [31:0] Register_inst226;
  reg [31:0] Register_inst227;
  reg [31:0] Register_inst228;
  reg [31:0] Register_inst229;
  reg [31:0] Register_inst230;
  reg [31:0] Register_inst231;
  reg [31:0] Register_inst232;
  reg [31:0] Register_inst233;
  reg [31:0] Register_inst234;
  reg [31:0] Register_inst235;
  reg [31:0] Register_inst236;
  reg [31:0] Register_inst237;
  reg [31:0] Register_inst238;
  reg [31:0] Register_inst239;
  reg [31:0] Register_inst240;
  reg [31:0] Register_inst241;
  reg [31:0] Register_inst242;
  reg [31:0] Register_inst243;
  reg [31:0] Register_inst244;
  reg [31:0] Register_inst245;
  reg [31:0] Register_inst246;
  reg [31:0] Register_inst247;
  reg [31:0] Register_inst248;
  reg [31:0] Register_inst249;
  reg [31:0] Register_inst250;
  reg [31:0] Register_inst251;
  reg [31:0] Register_inst252;
  reg [31:0] Register_inst253;
  reg [31:0] Register_inst254;
  reg [31:0] Register_inst255;

  always_ff @(posedge CLK or posedge ASYNCRESET) begin
    if (ASYNCRESET) begin
      Register_inst0 <= 32'h0;
      Register_inst1 <= 32'h0;
      Register_inst2 <= 32'h0;
      Register_inst3 <= 32'h0;
      Register_inst4 <= 32'h0;
      Register_inst5 <= 32'h0;
      Register_inst6 <= 32'h0;
      Register_inst7 <= 32'h0;
      Register_inst8 <= 32'h0;
      Register_inst9 <= 32'h0;
      Register_inst10 <= 32'h0;
      Register_inst11 <= 32'h0;
      Register_inst12 <= 32'h0;
      Register_inst13 <= 32'h0;
      Register_inst14 <= 32'h0;
      Register_inst15 <= 32'h0;
      Register_inst16 <= 32'h0;
      Register_inst17 <= 32'h0;
      Register_inst18 <= 32'h0;
      Register_inst19 <= 32'h0;
      Register_inst20 <= 32'h0;
      Register_inst21 <= 32'h0;
      Register_inst22 <= 32'h0;
      Register_inst23 <= 32'h0;
      Register_inst24 <= 32'h0;
      Register_inst25 <= 32'h0;
      Register_inst26 <= 32'h0;
      Register_inst27 <= 32'h0;
      Register_inst28 <= 32'h0;
      Register_inst29 <= 32'h0;
      Register_inst30 <= 32'h0;
      Register_inst31 <= 32'h0;
      Register_inst32 <= 32'h0;
      Register_inst33 <= 32'h0;
      Register_inst34 <= 32'h0;
      Register_inst35 <= 32'h0;
      Register_inst36 <= 32'h0;
      Register_inst37 <= 32'h0;
      Register_inst38 <= 32'h0;
      Register_inst39 <= 32'h0;
      Register_inst40 <= 32'h0;
      Register_inst41 <= 32'h0;
      Register_inst42 <= 32'h0;
      Register_inst43 <= 32'h0;
      Register_inst44 <= 32'h0;
      Register_inst45 <= 32'h0;
      Register_inst46 <= 32'h0;
      Register_inst47 <= 32'h0;
      Register_inst48 <= 32'h0;
      Register_inst49 <= 32'h0;
      Register_inst50 <= 32'h0;
      Register_inst51 <= 32'h0;
      Register_inst52 <= 32'h0;
      Register_inst53 <= 32'h0;
      Register_inst54 <= 32'h0;
      Register_inst55 <= 32'h0;
      Register_inst56 <= 32'h0;
      Register_inst57 <= 32'h0;
      Register_inst58 <= 32'h0;
      Register_inst59 <= 32'h0;
      Register_inst60 <= 32'h0;
      Register_inst61 <= 32'h0;
      Register_inst62 <= 32'h0;
      Register_inst63 <= 32'h0;
      Register_inst64 <= 32'h0;
      Register_inst65 <= 32'h0;
      Register_inst66 <= 32'h0;
      Register_inst67 <= 32'h0;
      Register_inst68 <= 32'h0;
      Register_inst69 <= 32'h0;
      Register_inst70 <= 32'h0;
      Register_inst71 <= 32'h0;
      Register_inst72 <= 32'h0;
      Register_inst73 <= 32'h0;
      Register_inst74 <= 32'h0;
      Register_inst75 <= 32'h0;
      Register_inst76 <= 32'h0;
      Register_inst77 <= 32'h0;
      Register_inst78 <= 32'h0;
      Register_inst79 <= 32'h0;
      Register_inst80 <= 32'h0;
      Register_inst81 <= 32'h0;
      Register_inst82 <= 32'h0;
      Register_inst83 <= 32'h0;
      Register_inst84 <= 32'h0;
      Register_inst85 <= 32'h0;
      Register_inst86 <= 32'h0;
      Register_inst87 <= 32'h0;
      Register_inst88 <= 32'h0;
      Register_inst89 <= 32'h0;
      Register_inst90 <= 32'h0;
      Register_inst91 <= 32'h0;
      Register_inst92 <= 32'h0;
      Register_inst93 <= 32'h0;
      Register_inst94 <= 32'h0;
      Register_inst95 <= 32'h0;
      Register_inst96 <= 32'h0;
      Register_inst97 <= 32'h0;
      Register_inst98 <= 32'h0;
      Register_inst99 <= 32'h0;
      Register_inst100 <= 32'h0;
      Register_inst101 <= 32'h0;
      Register_inst102 <= 32'h0;
      Register_inst103 <= 32'h0;
      Register_inst104 <= 32'h0;
      Register_inst105 <= 32'h0;
      Register_inst106 <= 32'h0;
      Register_inst107 <= 32'h0;
      Register_inst108 <= 32'h0;
      Register_inst109 <= 32'h0;
      Register_inst110 <= 32'h0;
      Register_inst111 <= 32'h0;
      Register_inst112 <= 32'h0;
      Register_inst113 <= 32'h0;
      Register_inst114 <= 32'h0;
      Register_inst115 <= 32'h0;
      Register_inst116 <= 32'h0;
      Register_inst117 <= 32'h0;
      Register_inst118 <= 32'h0;
      Register_inst119 <= 32'h0;
      Register_inst120 <= 32'h0;
      Register_inst121 <= 32'h0;
      Register_inst122 <= 32'h0;
      Register_inst123 <= 32'h0;
      Register_inst124 <= 32'h0;
      Register_inst125 <= 32'h0;
      Register_inst126 <= 32'h0;
      Register_inst127 <= 32'h0;
      Register_inst128 <= 32'h0;
      Register_inst129 <= 32'h0;
      Register_inst130 <= 32'h0;
      Register_inst131 <= 32'h0;
      Register_inst132 <= 32'h0;
      Register_inst133 <= 32'h0;
      Register_inst134 <= 32'h0;
      Register_inst135 <= 32'h0;
      Register_inst136 <= 32'h0;
      Register_inst137 <= 32'h0;
      Register_inst138 <= 32'h0;
      Register_inst139 <= 32'h0;
      Register_inst140 <= 32'h0;
      Register_inst141 <= 32'h0;
      Register_inst142 <= 32'h0;
      Register_inst143 <= 32'h0;
      Register_inst144 <= 32'h0;
      Register_inst145 <= 32'h0;
      Register_inst146 <= 32'h0;
      Register_inst147 <= 32'h0;
      Register_inst148 <= 32'h0;
      Register_inst149 <= 32'h0;
      Register_inst150 <= 32'h0;
      Register_inst151 <= 32'h0;
      Register_inst152 <= 32'h0;
      Register_inst153 <= 32'h0;
      Register_inst154 <= 32'h0;
      Register_inst155 <= 32'h0;
      Register_inst156 <= 32'h0;
      Register_inst157 <= 32'h0;
      Register_inst158 <= 32'h0;
      Register_inst159 <= 32'h0;
      Register_inst160 <= 32'h0;
      Register_inst161 <= 32'h0;
      Register_inst162 <= 32'h0;
      Register_inst163 <= 32'h0;
      Register_inst164 <= 32'h0;
      Register_inst165 <= 32'h0;
      Register_inst166 <= 32'h0;
      Register_inst167 <= 32'h0;
      Register_inst168 <= 32'h0;
      Register_inst169 <= 32'h0;
      Register_inst170 <= 32'h0;
      Register_inst171 <= 32'h0;
      Register_inst172 <= 32'h0;
      Register_inst173 <= 32'h0;
      Register_inst174 <= 32'h0;
      Register_inst175 <= 32'h0;
      Register_inst176 <= 32'h0;
      Register_inst177 <= 32'h0;
      Register_inst178 <= 32'h0;
      Register_inst179 <= 32'h0;
      Register_inst180 <= 32'h0;
      Register_inst181 <= 32'h0;
      Register_inst182 <= 32'h0;
      Register_inst183 <= 32'h0;
      Register_inst184 <= 32'h0;
      Register_inst185 <= 32'h0;
      Register_inst186 <= 32'h0;
      Register_inst187 <= 32'h0;
      Register_inst188 <= 32'h0;
      Register_inst189 <= 32'h0;
      Register_inst190 <= 32'h0;
      Register_inst191 <= 32'h0;
      Register_inst192 <= 32'h0;
      Register_inst193 <= 32'h0;
      Register_inst194 <= 32'h0;
      Register_inst195 <= 32'h0;
      Register_inst196 <= 32'h0;
      Register_inst197 <= 32'h0;
      Register_inst198 <= 32'h0;
      Register_inst199 <= 32'h0;
      Register_inst200 <= 32'h0;
      Register_inst201 <= 32'h0;
      Register_inst202 <= 32'h0;
      Register_inst203 <= 32'h0;
      Register_inst204 <= 32'h0;
      Register_inst205 <= 32'h0;
      Register_inst206 <= 32'h0;
      Register_inst207 <= 32'h0;
      Register_inst208 <= 32'h0;
      Register_inst209 <= 32'h0;
      Register_inst210 <= 32'h0;
      Register_inst211 <= 32'h0;
      Register_inst212 <= 32'h0;
      Register_inst213 <= 32'h0;
      Register_inst214 <= 32'h0;
      Register_inst215 <= 32'h0;
      Register_inst216 <= 32'h0;
      Register_inst217 <= 32'h0;
      Register_inst218 <= 32'h0;
      Register_inst219 <= 32'h0;
      Register_inst220 <= 32'h0;
      Register_inst221 <= 32'h0;
      Register_inst222 <= 32'h0;
      Register_inst223 <= 32'h0;
      Register_inst224 <= 32'h0;
      Register_inst225 <= 32'h0;
      Register_inst226 <= 32'h0;
      Register_inst227 <= 32'h0;
      Register_inst228 <= 32'h0;
      Register_inst229 <= 32'h0;
      Register_inst230 <= 32'h0;
      Register_inst231 <= 32'h0;
      Register_inst232 <= 32'h0;
      Register_inst233 <= 32'h0;
      Register_inst234 <= 32'h0;
      Register_inst235 <= 32'h0;
      Register_inst236 <= 32'h0;
      Register_inst237 <= 32'h0;
      Register_inst238 <= 32'h0;
      Register_inst239 <= 32'h0;
      Register_inst240 <= 32'h0;
      Register_inst241 <= 32'h0;
      Register_inst242 <= 32'h0;
      Register_inst243 <= 32'h0;
      Register_inst244 <= 32'h0;
      Register_inst245 <= 32'h0;
      Register_inst246 <= 32'h0;
      Register_inst247 <= 32'h0;
      Register_inst248 <= 32'h0;
      Register_inst249 <= 32'h0;
      Register_inst250 <= 32'h0;
      Register_inst251 <= 32'h0;
      Register_inst252 <= 32'h0;
      Register_inst253 <= 32'h0;
      Register_inst254 <= 32'h0;
      Register_inst255 <= 32'h0;
    end
    else begin
      automatic logic [31:0]      _T_1 = write_0.data;
      automatic logic [7:0]       _T_2 = write_0.addr;
      automatic logic [1:0][31:0] _T_3 = {{Register_inst0}, {_T_1}};
      automatic logic [1:0][31:0] _T_4 = {{Register_inst1}, {_T_1}};
      automatic logic [1:0][31:0] _T_5 = {{Register_inst2}, {_T_1}};
      automatic logic [1:0][31:0] _T_6 = {{Register_inst3}, {_T_1}};
      automatic logic [1:0][31:0] _T_7 = {{Register_inst4}, {_T_1}};
      automatic logic [1:0][31:0] _T_8 = {{Register_inst5}, {_T_1}};
      automatic logic [1:0][31:0] _T_9 = {{Register_inst6}, {_T_1}};
      automatic logic [1:0][31:0] _T_10 = {{Register_inst7}, {_T_1}};
      automatic logic [1:0][31:0] _T_11 = {{Register_inst8}, {_T_1}};
      automatic logic [1:0][31:0] _T_12 = {{Register_inst9}, {_T_1}};
      automatic logic [1:0][31:0] _T_13 = {{Register_inst10}, {_T_1}};
      automatic logic [1:0][31:0] _T_14 = {{Register_inst11}, {_T_1}};
      automatic logic [1:0][31:0] _T_15 = {{Register_inst12}, {_T_1}};
      automatic logic [1:0][31:0] _T_16 = {{Register_inst13}, {_T_1}};
      automatic logic [1:0][31:0] _T_17 = {{Register_inst14}, {_T_1}};
      automatic logic [1:0][31:0] _T_18 = {{Register_inst15}, {_T_1}};
      automatic logic [1:0][31:0] _T_19 = {{Register_inst16}, {_T_1}};
      automatic logic [1:0][31:0] _T_20 = {{Register_inst17}, {_T_1}};
      automatic logic [1:0][31:0] _T_21 = {{Register_inst18}, {_T_1}};
      automatic logic [1:0][31:0] _T_22 = {{Register_inst19}, {_T_1}};
      automatic logic [1:0][31:0] _T_23 = {{Register_inst20}, {_T_1}};
      automatic logic [1:0][31:0] _T_24 = {{Register_inst21}, {_T_1}};
      automatic logic [1:0][31:0] _T_25 = {{Register_inst22}, {_T_1}};
      automatic logic [1:0][31:0] _T_26 = {{Register_inst23}, {_T_1}};
      automatic logic [1:0][31:0] _T_27 = {{Register_inst24}, {_T_1}};
      automatic logic [1:0][31:0] _T_28 = {{Register_inst25}, {_T_1}};
      automatic logic [1:0][31:0] _T_29 = {{Register_inst26}, {_T_1}};
      automatic logic [1:0][31:0] _T_30 = {{Register_inst27}, {_T_1}};
      automatic logic [1:0][31:0] _T_31 = {{Register_inst28}, {_T_1}};
      automatic logic [1:0][31:0] _T_32 = {{Register_inst29}, {_T_1}};
      automatic logic [1:0][31:0] _T_33 = {{Register_inst30}, {_T_1}};
      automatic logic [1:0][31:0] _T_34 = {{Register_inst31}, {_T_1}};
      automatic logic [1:0][31:0] _T_35 = {{Register_inst32}, {_T_1}};
      automatic logic [1:0][31:0] _T_36 = {{Register_inst33}, {_T_1}};
      automatic logic [1:0][31:0] _T_37 = {{Register_inst34}, {_T_1}};
      automatic logic [1:0][31:0] _T_38 = {{Register_inst35}, {_T_1}};
      automatic logic [1:0][31:0] _T_39 = {{Register_inst36}, {_T_1}};
      automatic logic [1:0][31:0] _T_40 = {{Register_inst37}, {_T_1}};
      automatic logic [1:0][31:0] _T_41 = {{Register_inst38}, {_T_1}};
      automatic logic [1:0][31:0] _T_42 = {{Register_inst39}, {_T_1}};
      automatic logic [1:0][31:0] _T_43 = {{Register_inst40}, {_T_1}};
      automatic logic [1:0][31:0] _T_44 = {{Register_inst41}, {_T_1}};
      automatic logic [1:0][31:0] _T_45 = {{Register_inst42}, {_T_1}};
      automatic logic [1:0][31:0] _T_46 = {{Register_inst43}, {_T_1}};
      automatic logic [1:0][31:0] _T_47 = {{Register_inst44}, {_T_1}};
      automatic logic [1:0][31:0] _T_48 = {{Register_inst45}, {_T_1}};
      automatic logic [1:0][31:0] _T_49 = {{Register_inst46}, {_T_1}};
      automatic logic [1:0][31:0] _T_50 = {{Register_inst47}, {_T_1}};
      automatic logic [1:0][31:0] _T_51 = {{Register_inst48}, {_T_1}};
      automatic logic [1:0][31:0] _T_52 = {{Register_inst49}, {_T_1}};
      automatic logic [1:0][31:0] _T_53 = {{Register_inst50}, {_T_1}};
      automatic logic [1:0][31:0] _T_54 = {{Register_inst51}, {_T_1}};
      automatic logic [1:0][31:0] _T_55 = {{Register_inst52}, {_T_1}};
      automatic logic [1:0][31:0] _T_56 = {{Register_inst53}, {_T_1}};
      automatic logic [1:0][31:0] _T_57 = {{Register_inst54}, {_T_1}};
      automatic logic [1:0][31:0] _T_58 = {{Register_inst55}, {_T_1}};
      automatic logic [1:0][31:0] _T_59 = {{Register_inst56}, {_T_1}};
      automatic logic [1:0][31:0] _T_60 = {{Register_inst57}, {_T_1}};
      automatic logic [1:0][31:0] _T_61 = {{Register_inst58}, {_T_1}};
      automatic logic [1:0][31:0] _T_62 = {{Register_inst59}, {_T_1}};
      automatic logic [1:0][31:0] _T_63 = {{Register_inst60}, {_T_1}};
      automatic logic [1:0][31:0] _T_64 = {{Register_inst61}, {_T_1}};
      automatic logic [1:0][31:0] _T_65 = {{Register_inst62}, {_T_1}};
      automatic logic [1:0][31:0] _T_66 = {{Register_inst63}, {_T_1}};
      automatic logic [1:0][31:0] _T_67 = {{Register_inst64}, {_T_1}};
      automatic logic [1:0][31:0] _T_68 = {{Register_inst65}, {_T_1}};
      automatic logic [1:0][31:0] _T_69 = {{Register_inst66}, {_T_1}};
      automatic logic [1:0][31:0] _T_70 = {{Register_inst67}, {_T_1}};
      automatic logic [1:0][31:0] _T_71 = {{Register_inst68}, {_T_1}};
      automatic logic [1:0][31:0] _T_72 = {{Register_inst69}, {_T_1}};
      automatic logic [1:0][31:0] _T_73 = {{Register_inst70}, {_T_1}};
      automatic logic [1:0][31:0] _T_74 = {{Register_inst71}, {_T_1}};
      automatic logic [1:0][31:0] _T_75 = {{Register_inst72}, {_T_1}};
      automatic logic [1:0][31:0] _T_76 = {{Register_inst73}, {_T_1}};
      automatic logic [1:0][31:0] _T_77 = {{Register_inst74}, {_T_1}};
      automatic logic [1:0][31:0] _T_78 = {{Register_inst75}, {_T_1}};
      automatic logic [1:0][31:0] _T_79 = {{Register_inst76}, {_T_1}};
      automatic logic [1:0][31:0] _T_80 = {{Register_inst77}, {_T_1}};
      automatic logic [1:0][31:0] _T_81 = {{Register_inst78}, {_T_1}};
      automatic logic [1:0][31:0] _T_82 = {{Register_inst79}, {_T_1}};
      automatic logic [1:0][31:0] _T_83 = {{Register_inst80}, {_T_1}};
      automatic logic [1:0][31:0] _T_84 = {{Register_inst81}, {_T_1}};
      automatic logic [1:0][31:0] _T_85 = {{Register_inst82}, {_T_1}};
      automatic logic [1:0][31:0] _T_86 = {{Register_inst83}, {_T_1}};
      automatic logic [1:0][31:0] _T_87 = {{Register_inst84}, {_T_1}};
      automatic logic [1:0][31:0] _T_88 = {{Register_inst85}, {_T_1}};
      automatic logic [1:0][31:0] _T_89 = {{Register_inst86}, {_T_1}};
      automatic logic [1:0][31:0] _T_90 = {{Register_inst87}, {_T_1}};
      automatic logic [1:0][31:0] _T_91 = {{Register_inst88}, {_T_1}};
      automatic logic [1:0][31:0] _T_92 = {{Register_inst89}, {_T_1}};
      automatic logic [1:0][31:0] _T_93 = {{Register_inst90}, {_T_1}};
      automatic logic [1:0][31:0] _T_94 = {{Register_inst91}, {_T_1}};
      automatic logic [1:0][31:0] _T_95 = {{Register_inst92}, {_T_1}};
      automatic logic [1:0][31:0] _T_96 = {{Register_inst93}, {_T_1}};
      automatic logic [1:0][31:0] _T_97 = {{Register_inst94}, {_T_1}};
      automatic logic [1:0][31:0] _T_98 = {{Register_inst95}, {_T_1}};
      automatic logic [1:0][31:0] _T_99 = {{Register_inst96}, {_T_1}};
      automatic logic [1:0][31:0] _T_100 = {{Register_inst97}, {_T_1}};
      automatic logic [1:0][31:0] _T_101 = {{Register_inst98}, {_T_1}};
      automatic logic [1:0][31:0] _T_102 = {{Register_inst99}, {_T_1}};
      automatic logic [1:0][31:0] _T_103 = {{Register_inst100}, {_T_1}};
      automatic logic [1:0][31:0] _T_104 = {{Register_inst101}, {_T_1}};
      automatic logic [1:0][31:0] _T_105 = {{Register_inst102}, {_T_1}};
      automatic logic [1:0][31:0] _T_106 = {{Register_inst103}, {_T_1}};
      automatic logic [1:0][31:0] _T_107 = {{Register_inst104}, {_T_1}};
      automatic logic [1:0][31:0] _T_108 = {{Register_inst105}, {_T_1}};
      automatic logic [1:0][31:0] _T_109 = {{Register_inst106}, {_T_1}};
      automatic logic [1:0][31:0] _T_110 = {{Register_inst107}, {_T_1}};
      automatic logic [1:0][31:0] _T_111 = {{Register_inst108}, {_T_1}};
      automatic logic [1:0][31:0] _T_112 = {{Register_inst109}, {_T_1}};
      automatic logic [1:0][31:0] _T_113 = {{Register_inst110}, {_T_1}};
      automatic logic [1:0][31:0] _T_114 = {{Register_inst111}, {_T_1}};
      automatic logic [1:0][31:0] _T_115 = {{Register_inst112}, {_T_1}};
      automatic logic [1:0][31:0] _T_116 = {{Register_inst113}, {_T_1}};
      automatic logic [1:0][31:0] _T_117 = {{Register_inst114}, {_T_1}};
      automatic logic [1:0][31:0] _T_118 = {{Register_inst115}, {_T_1}};
      automatic logic [1:0][31:0] _T_119 = {{Register_inst116}, {_T_1}};
      automatic logic [1:0][31:0] _T_120 = {{Register_inst117}, {_T_1}};
      automatic logic [1:0][31:0] _T_121 = {{Register_inst118}, {_T_1}};
      automatic logic [1:0][31:0] _T_122 = {{Register_inst119}, {_T_1}};
      automatic logic [1:0][31:0] _T_123 = {{Register_inst120}, {_T_1}};
      automatic logic [1:0][31:0] _T_124 = {{Register_inst121}, {_T_1}};
      automatic logic [1:0][31:0] _T_125 = {{Register_inst122}, {_T_1}};
      automatic logic [1:0][31:0] _T_126 = {{Register_inst123}, {_T_1}};
      automatic logic [1:0][31:0] _T_127 = {{Register_inst124}, {_T_1}};
      automatic logic [1:0][31:0] _T_128 = {{Register_inst125}, {_T_1}};
      automatic logic [1:0][31:0] _T_129 = {{Register_inst126}, {_T_1}};
      automatic logic [1:0][31:0] _T_130 = {{Register_inst127}, {_T_1}};
      automatic logic [1:0][31:0] _T_131 = {{Register_inst128}, {_T_1}};
      automatic logic [1:0][31:0] _T_132 = {{Register_inst129}, {_T_1}};
      automatic logic [1:0][31:0] _T_133 = {{Register_inst130}, {_T_1}};
      automatic logic [1:0][31:0] _T_134 = {{Register_inst131}, {_T_1}};
      automatic logic [1:0][31:0] _T_135 = {{Register_inst132}, {_T_1}};
      automatic logic [1:0][31:0] _T_136 = {{Register_inst133}, {_T_1}};
      automatic logic [1:0][31:0] _T_137 = {{Register_inst134}, {_T_1}};
      automatic logic [1:0][31:0] _T_138 = {{Register_inst135}, {_T_1}};
      automatic logic [1:0][31:0] _T_139 = {{Register_inst136}, {_T_1}};
      automatic logic [1:0][31:0] _T_140 = {{Register_inst137}, {_T_1}};
      automatic logic [1:0][31:0] _T_141 = {{Register_inst138}, {_T_1}};
      automatic logic [1:0][31:0] _T_142 = {{Register_inst139}, {_T_1}};
      automatic logic [1:0][31:0] _T_143 = {{Register_inst140}, {_T_1}};
      automatic logic [1:0][31:0] _T_144 = {{Register_inst141}, {_T_1}};
      automatic logic [1:0][31:0] _T_145 = {{Register_inst142}, {_T_1}};
      automatic logic [1:0][31:0] _T_146 = {{Register_inst143}, {_T_1}};
      automatic logic [1:0][31:0] _T_147 = {{Register_inst144}, {_T_1}};
      automatic logic [1:0][31:0] _T_148 = {{Register_inst145}, {_T_1}};
      automatic logic [1:0][31:0] _T_149 = {{Register_inst146}, {_T_1}};
      automatic logic [1:0][31:0] _T_150 = {{Register_inst147}, {_T_1}};
      automatic logic [1:0][31:0] _T_151 = {{Register_inst148}, {_T_1}};
      automatic logic [1:0][31:0] _T_152 = {{Register_inst149}, {_T_1}};
      automatic logic [1:0][31:0] _T_153 = {{Register_inst150}, {_T_1}};
      automatic logic [1:0][31:0] _T_154 = {{Register_inst151}, {_T_1}};
      automatic logic [1:0][31:0] _T_155 = {{Register_inst152}, {_T_1}};
      automatic logic [1:0][31:0] _T_156 = {{Register_inst153}, {_T_1}};
      automatic logic [1:0][31:0] _T_157 = {{Register_inst154}, {_T_1}};
      automatic logic [1:0][31:0] _T_158 = {{Register_inst155}, {_T_1}};
      automatic logic [1:0][31:0] _T_159 = {{Register_inst156}, {_T_1}};
      automatic logic [1:0][31:0] _T_160 = {{Register_inst157}, {_T_1}};
      automatic logic [1:0][31:0] _T_161 = {{Register_inst158}, {_T_1}};
      automatic logic [1:0][31:0] _T_162 = {{Register_inst159}, {_T_1}};
      automatic logic [1:0][31:0] _T_163 = {{Register_inst160}, {_T_1}};
      automatic logic [1:0][31:0] _T_164 = {{Register_inst161}, {_T_1}};
      automatic logic [1:0][31:0] _T_165 = {{Register_inst162}, {_T_1}};
      automatic logic [1:0][31:0] _T_166 = {{Register_inst163}, {_T_1}};
      automatic logic [1:0][31:0] _T_167 = {{Register_inst164}, {_T_1}};
      automatic logic [1:0][31:0] _T_168 = {{Register_inst165}, {_T_1}};
      automatic logic [1:0][31:0] _T_169 = {{Register_inst166}, {_T_1}};
      automatic logic [1:0][31:0] _T_170 = {{Register_inst167}, {_T_1}};
      automatic logic [1:0][31:0] _T_171 = {{Register_inst168}, {_T_1}};
      automatic logic [1:0][31:0] _T_172 = {{Register_inst169}, {_T_1}};
      automatic logic [1:0][31:0] _T_173 = {{Register_inst170}, {_T_1}};
      automatic logic [1:0][31:0] _T_174 = {{Register_inst171}, {_T_1}};
      automatic logic [1:0][31:0] _T_175 = {{Register_inst172}, {_T_1}};
      automatic logic [1:0][31:0] _T_176 = {{Register_inst173}, {_T_1}};
      automatic logic [1:0][31:0] _T_177 = {{Register_inst174}, {_T_1}};
      automatic logic [1:0][31:0] _T_178 = {{Register_inst175}, {_T_1}};
      automatic logic [1:0][31:0] _T_179 = {{Register_inst176}, {_T_1}};
      automatic logic [1:0][31:0] _T_180 = {{Register_inst177}, {_T_1}};
      automatic logic [1:0][31:0] _T_181 = {{Register_inst178}, {_T_1}};
      automatic logic [1:0][31:0] _T_182 = {{Register_inst179}, {_T_1}};
      automatic logic [1:0][31:0] _T_183 = {{Register_inst180}, {_T_1}};
      automatic logic [1:0][31:0] _T_184 = {{Register_inst181}, {_T_1}};
      automatic logic [1:0][31:0] _T_185 = {{Register_inst182}, {_T_1}};
      automatic logic [1:0][31:0] _T_186 = {{Register_inst183}, {_T_1}};
      automatic logic [1:0][31:0] _T_187 = {{Register_inst184}, {_T_1}};
      automatic logic [1:0][31:0] _T_188 = {{Register_inst185}, {_T_1}};
      automatic logic [1:0][31:0] _T_189 = {{Register_inst186}, {_T_1}};
      automatic logic [1:0][31:0] _T_190 = {{Register_inst187}, {_T_1}};
      automatic logic [1:0][31:0] _T_191 = {{Register_inst188}, {_T_1}};
      automatic logic [1:0][31:0] _T_192 = {{Register_inst189}, {_T_1}};
      automatic logic [1:0][31:0] _T_193 = {{Register_inst190}, {_T_1}};
      automatic logic [1:0][31:0] _T_194 = {{Register_inst191}, {_T_1}};
      automatic logic [1:0][31:0] _T_195 = {{Register_inst192}, {_T_1}};
      automatic logic [1:0][31:0] _T_196 = {{Register_inst193}, {_T_1}};
      automatic logic [1:0][31:0] _T_197 = {{Register_inst194}, {_T_1}};
      automatic logic [1:0][31:0] _T_198 = {{Register_inst195}, {_T_1}};
      automatic logic [1:0][31:0] _T_199 = {{Register_inst196}, {_T_1}};
      automatic logic [1:0][31:0] _T_200 = {{Register_inst197}, {_T_1}};
      automatic logic [1:0][31:0] _T_201 = {{Register_inst198}, {_T_1}};
      automatic logic [1:0][31:0] _T_202 = {{Register_inst199}, {_T_1}};
      automatic logic [1:0][31:0] _T_203 = {{Register_inst200}, {_T_1}};
      automatic logic [1:0][31:0] _T_204 = {{Register_inst201}, {_T_1}};
      automatic logic [1:0][31:0] _T_205 = {{Register_inst202}, {_T_1}};
      automatic logic [1:0][31:0] _T_206 = {{Register_inst203}, {_T_1}};
      automatic logic [1:0][31:0] _T_207 = {{Register_inst204}, {_T_1}};
      automatic logic [1:0][31:0] _T_208 = {{Register_inst205}, {_T_1}};
      automatic logic [1:0][31:0] _T_209 = {{Register_inst206}, {_T_1}};
      automatic logic [1:0][31:0] _T_210 = {{Register_inst207}, {_T_1}};
      automatic logic [1:0][31:0] _T_211 = {{Register_inst208}, {_T_1}};
      automatic logic [1:0][31:0] _T_212 = {{Register_inst209}, {_T_1}};
      automatic logic [1:0][31:0] _T_213 = {{Register_inst210}, {_T_1}};
      automatic logic [1:0][31:0] _T_214 = {{Register_inst211}, {_T_1}};
      automatic logic [1:0][31:0] _T_215 = {{Register_inst212}, {_T_1}};
      automatic logic [1:0][31:0] _T_216 = {{Register_inst213}, {_T_1}};
      automatic logic [1:0][31:0] _T_217 = {{Register_inst214}, {_T_1}};
      automatic logic [1:0][31:0] _T_218 = {{Register_inst215}, {_T_1}};
      automatic logic [1:0][31:0] _T_219 = {{Register_inst216}, {_T_1}};
      automatic logic [1:0][31:0] _T_220 = {{Register_inst217}, {_T_1}};
      automatic logic [1:0][31:0] _T_221 = {{Register_inst218}, {_T_1}};
      automatic logic [1:0][31:0] _T_222 = {{Register_inst219}, {_T_1}};
      automatic logic [1:0][31:0] _T_223 = {{Register_inst220}, {_T_1}};
      automatic logic [1:0][31:0] _T_224 = {{Register_inst221}, {_T_1}};
      automatic logic [1:0][31:0] _T_225 = {{Register_inst222}, {_T_1}};
      automatic logic [1:0][31:0] _T_226 = {{Register_inst223}, {_T_1}};
      automatic logic [1:0][31:0] _T_227 = {{Register_inst224}, {_T_1}};
      automatic logic [1:0][31:0] _T_228 = {{Register_inst225}, {_T_1}};
      automatic logic [1:0][31:0] _T_229 = {{Register_inst226}, {_T_1}};
      automatic logic [1:0][31:0] _T_230 = {{Register_inst227}, {_T_1}};
      automatic logic [1:0][31:0] _T_231 = {{Register_inst228}, {_T_1}};
      automatic logic [1:0][31:0] _T_232 = {{Register_inst229}, {_T_1}};
      automatic logic [1:0][31:0] _T_233 = {{Register_inst230}, {_T_1}};
      automatic logic [1:0][31:0] _T_234 = {{Register_inst231}, {_T_1}};
      automatic logic [1:0][31:0] _T_235 = {{Register_inst232}, {_T_1}};
      automatic logic [1:0][31:0] _T_236 = {{Register_inst233}, {_T_1}};
      automatic logic [1:0][31:0] _T_237 = {{Register_inst234}, {_T_1}};
      automatic logic [1:0][31:0] _T_238 = {{Register_inst235}, {_T_1}};
      automatic logic [1:0][31:0] _T_239 = {{Register_inst236}, {_T_1}};
      automatic logic [1:0][31:0] _T_240 = {{Register_inst237}, {_T_1}};
      automatic logic [1:0][31:0] _T_241 = {{Register_inst238}, {_T_1}};
      automatic logic [1:0][31:0] _T_242 = {{Register_inst239}, {_T_1}};
      automatic logic [1:0][31:0] _T_243 = {{Register_inst240}, {_T_1}};
      automatic logic [1:0][31:0] _T_244 = {{Register_inst241}, {_T_1}};
      automatic logic [1:0][31:0] _T_245 = {{Register_inst242}, {_T_1}};
      automatic logic [1:0][31:0] _T_246 = {{Register_inst243}, {_T_1}};
      automatic logic [1:0][31:0] _T_247 = {{Register_inst244}, {_T_1}};
      automatic logic [1:0][31:0] _T_248 = {{Register_inst245}, {_T_1}};
      automatic logic [1:0][31:0] _T_249 = {{Register_inst246}, {_T_1}};
      automatic logic [1:0][31:0] _T_250 = {{Register_inst247}, {_T_1}};
      automatic logic [1:0][31:0] _T_251 = {{Register_inst248}, {_T_1}};
      automatic logic [1:0][31:0] _T_252 = {{Register_inst249}, {_T_1}};
      automatic logic [1:0][31:0] _T_253 = {{Register_inst250}, {_T_1}};
      automatic logic [1:0][31:0] _T_254 = {{Register_inst251}, {_T_1}};
      automatic logic [1:0][31:0] _T_255 = {{Register_inst252}, {_T_1}};
      automatic logic [1:0][31:0] _T_256 = {{Register_inst253}, {_T_1}};
      automatic logic [1:0][31:0] _T_257 = {{Register_inst254}, {_T_1}};
      automatic logic [1:0][31:0] _T_258 = {{Register_inst255}, {_T_1}};

      Register_inst0 <= _T_3[_T_2 == 8'h0 & write_0_en];
      Register_inst1 <= _T_4[_T_2 == 8'h1 & write_0_en];
      Register_inst2 <= _T_5[_T_2 == 8'h2 & write_0_en];
      Register_inst3 <= _T_6[_T_2 == 8'h3 & write_0_en];
      Register_inst4 <= _T_7[_T_2 == 8'h4 & write_0_en];
      Register_inst5 <= _T_8[_T_2 == 8'h5 & write_0_en];
      Register_inst6 <= _T_9[_T_2 == 8'h6 & write_0_en];
      Register_inst7 <= _T_10[_T_2 == 8'h7 & write_0_en];
      Register_inst8 <= _T_11[_T_2 == 8'h8 & write_0_en];
      Register_inst9 <= _T_12[_T_2 == 8'h9 & write_0_en];
      Register_inst10 <= _T_13[_T_2 == 8'hA & write_0_en];
      Register_inst11 <= _T_14[_T_2 == 8'hB & write_0_en];
      Register_inst12 <= _T_15[_T_2 == 8'hC & write_0_en];
      Register_inst13 <= _T_16[_T_2 == 8'hD & write_0_en];
      Register_inst14 <= _T_17[_T_2 == 8'hE & write_0_en];
      Register_inst15 <= _T_18[_T_2 == 8'hF & write_0_en];
      Register_inst16 <= _T_19[_T_2 == 8'h10 & write_0_en];
      Register_inst17 <= _T_20[_T_2 == 8'h11 & write_0_en];
      Register_inst18 <= _T_21[_T_2 == 8'h12 & write_0_en];
      Register_inst19 <= _T_22[_T_2 == 8'h13 & write_0_en];
      Register_inst20 <= _T_23[_T_2 == 8'h14 & write_0_en];
      Register_inst21 <= _T_24[_T_2 == 8'h15 & write_0_en];
      Register_inst22 <= _T_25[_T_2 == 8'h16 & write_0_en];
      Register_inst23 <= _T_26[_T_2 == 8'h17 & write_0_en];
      Register_inst24 <= _T_27[_T_2 == 8'h18 & write_0_en];
      Register_inst25 <= _T_28[_T_2 == 8'h19 & write_0_en];
      Register_inst26 <= _T_29[_T_2 == 8'h1A & write_0_en];
      Register_inst27 <= _T_30[_T_2 == 8'h1B & write_0_en];
      Register_inst28 <= _T_31[_T_2 == 8'h1C & write_0_en];
      Register_inst29 <= _T_32[_T_2 == 8'h1D & write_0_en];
      Register_inst30 <= _T_33[_T_2 == 8'h1E & write_0_en];
      Register_inst31 <= _T_34[_T_2 == 8'h1F & write_0_en];
      Register_inst32 <= _T_35[_T_2 == 8'h20 & write_0_en];
      Register_inst33 <= _T_36[_T_2 == 8'h21 & write_0_en];
      Register_inst34 <= _T_37[_T_2 == 8'h22 & write_0_en];
      Register_inst35 <= _T_38[_T_2 == 8'h23 & write_0_en];
      Register_inst36 <= _T_39[_T_2 == 8'h24 & write_0_en];
      Register_inst37 <= _T_40[_T_2 == 8'h25 & write_0_en];
      Register_inst38 <= _T_41[_T_2 == 8'h26 & write_0_en];
      Register_inst39 <= _T_42[_T_2 == 8'h27 & write_0_en];
      Register_inst40 <= _T_43[_T_2 == 8'h28 & write_0_en];
      Register_inst41 <= _T_44[_T_2 == 8'h29 & write_0_en];
      Register_inst42 <= _T_45[_T_2 == 8'h2A & write_0_en];
      Register_inst43 <= _T_46[_T_2 == 8'h2B & write_0_en];
      Register_inst44 <= _T_47[_T_2 == 8'h2C & write_0_en];
      Register_inst45 <= _T_48[_T_2 == 8'h2D & write_0_en];
      Register_inst46 <= _T_49[_T_2 == 8'h2E & write_0_en];
      Register_inst47 <= _T_50[_T_2 == 8'h2F & write_0_en];
      Register_inst48 <= _T_51[_T_2 == 8'h30 & write_0_en];
      Register_inst49 <= _T_52[_T_2 == 8'h31 & write_0_en];
      Register_inst50 <= _T_53[_T_2 == 8'h32 & write_0_en];
      Register_inst51 <= _T_54[_T_2 == 8'h33 & write_0_en];
      Register_inst52 <= _T_55[_T_2 == 8'h34 & write_0_en];
      Register_inst53 <= _T_56[_T_2 == 8'h35 & write_0_en];
      Register_inst54 <= _T_57[_T_2 == 8'h36 & write_0_en];
      Register_inst55 <= _T_58[_T_2 == 8'h37 & write_0_en];
      Register_inst56 <= _T_59[_T_2 == 8'h38 & write_0_en];
      Register_inst57 <= _T_60[_T_2 == 8'h39 & write_0_en];
      Register_inst58 <= _T_61[_T_2 == 8'h3A & write_0_en];
      Register_inst59 <= _T_62[_T_2 == 8'h3B & write_0_en];
      Register_inst60 <= _T_63[_T_2 == 8'h3C & write_0_en];
      Register_inst61 <= _T_64[_T_2 == 8'h3D & write_0_en];
      Register_inst62 <= _T_65[_T_2 == 8'h3E & write_0_en];
      Register_inst63 <= _T_66[_T_2 == 8'h3F & write_0_en];
      Register_inst64 <= _T_67[_T_2 == 8'h40 & write_0_en];
      Register_inst65 <= _T_68[_T_2 == 8'h41 & write_0_en];
      Register_inst66 <= _T_69[_T_2 == 8'h42 & write_0_en];
      Register_inst67 <= _T_70[_T_2 == 8'h43 & write_0_en];
      Register_inst68 <= _T_71[_T_2 == 8'h44 & write_0_en];
      Register_inst69 <= _T_72[_T_2 == 8'h45 & write_0_en];
      Register_inst70 <= _T_73[_T_2 == 8'h46 & write_0_en];
      Register_inst71 <= _T_74[_T_2 == 8'h47 & write_0_en];
      Register_inst72 <= _T_75[_T_2 == 8'h48 & write_0_en];
      Register_inst73 <= _T_76[_T_2 == 8'h49 & write_0_en];
      Register_inst74 <= _T_77[_T_2 == 8'h4A & write_0_en];
      Register_inst75 <= _T_78[_T_2 == 8'h4B & write_0_en];
      Register_inst76 <= _T_79[_T_2 == 8'h4C & write_0_en];
      Register_inst77 <= _T_80[_T_2 == 8'h4D & write_0_en];
      Register_inst78 <= _T_81[_T_2 == 8'h4E & write_0_en];
      Register_inst79 <= _T_82[_T_2 == 8'h4F & write_0_en];
      Register_inst80 <= _T_83[_T_2 == 8'h50 & write_0_en];
      Register_inst81 <= _T_84[_T_2 == 8'h51 & write_0_en];
      Register_inst82 <= _T_85[_T_2 == 8'h52 & write_0_en];
      Register_inst83 <= _T_86[_T_2 == 8'h53 & write_0_en];
      Register_inst84 <= _T_87[_T_2 == 8'h54 & write_0_en];
      Register_inst85 <= _T_88[_T_2 == 8'h55 & write_0_en];
      Register_inst86 <= _T_89[_T_2 == 8'h56 & write_0_en];
      Register_inst87 <= _T_90[_T_2 == 8'h57 & write_0_en];
      Register_inst88 <= _T_91[_T_2 == 8'h58 & write_0_en];
      Register_inst89 <= _T_92[_T_2 == 8'h59 & write_0_en];
      Register_inst90 <= _T_93[_T_2 == 8'h5A & write_0_en];
      Register_inst91 <= _T_94[_T_2 == 8'h5B & write_0_en];
      Register_inst92 <= _T_95[_T_2 == 8'h5C & write_0_en];
      Register_inst93 <= _T_96[_T_2 == 8'h5D & write_0_en];
      Register_inst94 <= _T_97[_T_2 == 8'h5E & write_0_en];
      Register_inst95 <= _T_98[_T_2 == 8'h5F & write_0_en];
      Register_inst96 <= _T_99[_T_2 == 8'h60 & write_0_en];
      Register_inst97 <= _T_100[_T_2 == 8'h61 & write_0_en];
      Register_inst98 <= _T_101[_T_2 == 8'h62 & write_0_en];
      Register_inst99 <= _T_102[_T_2 == 8'h63 & write_0_en];
      Register_inst100 <= _T_103[_T_2 == 8'h64 & write_0_en];
      Register_inst101 <= _T_104[_T_2 == 8'h65 & write_0_en];
      Register_inst102 <= _T_105[_T_2 == 8'h66 & write_0_en];
      Register_inst103 <= _T_106[_T_2 == 8'h67 & write_0_en];
      Register_inst104 <= _T_107[_T_2 == 8'h68 & write_0_en];
      Register_inst105 <= _T_108[_T_2 == 8'h69 & write_0_en];
      Register_inst106 <= _T_109[_T_2 == 8'h6A & write_0_en];
      Register_inst107 <= _T_110[_T_2 == 8'h6B & write_0_en];
      Register_inst108 <= _T_111[_T_2 == 8'h6C & write_0_en];
      Register_inst109 <= _T_112[_T_2 == 8'h6D & write_0_en];
      Register_inst110 <= _T_113[_T_2 == 8'h6E & write_0_en];
      Register_inst111 <= _T_114[_T_2 == 8'h6F & write_0_en];
      Register_inst112 <= _T_115[_T_2 == 8'h70 & write_0_en];
      Register_inst113 <= _T_116[_T_2 == 8'h71 & write_0_en];
      Register_inst114 <= _T_117[_T_2 == 8'h72 & write_0_en];
      Register_inst115 <= _T_118[_T_2 == 8'h73 & write_0_en];
      Register_inst116 <= _T_119[_T_2 == 8'h74 & write_0_en];
      Register_inst117 <= _T_120[_T_2 == 8'h75 & write_0_en];
      Register_inst118 <= _T_121[_T_2 == 8'h76 & write_0_en];
      Register_inst119 <= _T_122[_T_2 == 8'h77 & write_0_en];
      Register_inst120 <= _T_123[_T_2 == 8'h78 & write_0_en];
      Register_inst121 <= _T_124[_T_2 == 8'h79 & write_0_en];
      Register_inst122 <= _T_125[_T_2 == 8'h7A & write_0_en];
      Register_inst123 <= _T_126[_T_2 == 8'h7B & write_0_en];
      Register_inst124 <= _T_127[_T_2 == 8'h7C & write_0_en];
      Register_inst125 <= _T_128[_T_2 == 8'h7D & write_0_en];
      Register_inst126 <= _T_129[_T_2 == 8'h7E & write_0_en];
      Register_inst127 <= _T_130[_T_2 == 8'h7F & write_0_en];
      Register_inst128 <= _T_131[_T_2 == 8'h80 & write_0_en];
      Register_inst129 <= _T_132[_T_2 == 8'h81 & write_0_en];
      Register_inst130 <= _T_133[_T_2 == 8'h82 & write_0_en];
      Register_inst131 <= _T_134[_T_2 == 8'h83 & write_0_en];
      Register_inst132 <= _T_135[_T_2 == 8'h84 & write_0_en];
      Register_inst133 <= _T_136[_T_2 == 8'h85 & write_0_en];
      Register_inst134 <= _T_137[_T_2 == 8'h86 & write_0_en];
      Register_inst135 <= _T_138[_T_2 == 8'h87 & write_0_en];
      Register_inst136 <= _T_139[_T_2 == 8'h88 & write_0_en];
      Register_inst137 <= _T_140[_T_2 == 8'h89 & write_0_en];
      Register_inst138 <= _T_141[_T_2 == 8'h8A & write_0_en];
      Register_inst139 <= _T_142[_T_2 == 8'h8B & write_0_en];
      Register_inst140 <= _T_143[_T_2 == 8'h8C & write_0_en];
      Register_inst141 <= _T_144[_T_2 == 8'h8D & write_0_en];
      Register_inst142 <= _T_145[_T_2 == 8'h8E & write_0_en];
      Register_inst143 <= _T_146[_T_2 == 8'h8F & write_0_en];
      Register_inst144 <= _T_147[_T_2 == 8'h90 & write_0_en];
      Register_inst145 <= _T_148[_T_2 == 8'h91 & write_0_en];
      Register_inst146 <= _T_149[_T_2 == 8'h92 & write_0_en];
      Register_inst147 <= _T_150[_T_2 == 8'h93 & write_0_en];
      Register_inst148 <= _T_151[_T_2 == 8'h94 & write_0_en];
      Register_inst149 <= _T_152[_T_2 == 8'h95 & write_0_en];
      Register_inst150 <= _T_153[_T_2 == 8'h96 & write_0_en];
      Register_inst151 <= _T_154[_T_2 == 8'h97 & write_0_en];
      Register_inst152 <= _T_155[_T_2 == 8'h98 & write_0_en];
      Register_inst153 <= _T_156[_T_2 == 8'h99 & write_0_en];
      Register_inst154 <= _T_157[_T_2 == 8'h9A & write_0_en];
      Register_inst155 <= _T_158[_T_2 == 8'h9B & write_0_en];
      Register_inst156 <= _T_159[_T_2 == 8'h9C & write_0_en];
      Register_inst157 <= _T_160[_T_2 == 8'h9D & write_0_en];
      Register_inst158 <= _T_161[_T_2 == 8'h9E & write_0_en];
      Register_inst159 <= _T_162[_T_2 == 8'h9F & write_0_en];
      Register_inst160 <= _T_163[_T_2 == 8'hA0 & write_0_en];
      Register_inst161 <= _T_164[_T_2 == 8'hA1 & write_0_en];
      Register_inst162 <= _T_165[_T_2 == 8'hA2 & write_0_en];
      Register_inst163 <= _T_166[_T_2 == 8'hA3 & write_0_en];
      Register_inst164 <= _T_167[_T_2 == 8'hA4 & write_0_en];
      Register_inst165 <= _T_168[_T_2 == 8'hA5 & write_0_en];
      Register_inst166 <= _T_169[_T_2 == 8'hA6 & write_0_en];
      Register_inst167 <= _T_170[_T_2 == 8'hA7 & write_0_en];
      Register_inst168 <= _T_171[_T_2 == 8'hA8 & write_0_en];
      Register_inst169 <= _T_172[_T_2 == 8'hA9 & write_0_en];
      Register_inst170 <= _T_173[_T_2 == 8'hAA & write_0_en];
      Register_inst171 <= _T_174[_T_2 == 8'hAB & write_0_en];
      Register_inst172 <= _T_175[_T_2 == 8'hAC & write_0_en];
      Register_inst173 <= _T_176[_T_2 == 8'hAD & write_0_en];
      Register_inst174 <= _T_177[_T_2 == 8'hAE & write_0_en];
      Register_inst175 <= _T_178[_T_2 == 8'hAF & write_0_en];
      Register_inst176 <= _T_179[_T_2 == 8'hB0 & write_0_en];
      Register_inst177 <= _T_180[_T_2 == 8'hB1 & write_0_en];
      Register_inst178 <= _T_181[_T_2 == 8'hB2 & write_0_en];
      Register_inst179 <= _T_182[_T_2 == 8'hB3 & write_0_en];
      Register_inst180 <= _T_183[_T_2 == 8'hB4 & write_0_en];
      Register_inst181 <= _T_184[_T_2 == 8'hB5 & write_0_en];
      Register_inst182 <= _T_185[_T_2 == 8'hB6 & write_0_en];
      Register_inst183 <= _T_186[_T_2 == 8'hB7 & write_0_en];
      Register_inst184 <= _T_187[_T_2 == 8'hB8 & write_0_en];
      Register_inst185 <= _T_188[_T_2 == 8'hB9 & write_0_en];
      Register_inst186 <= _T_189[_T_2 == 8'hBA & write_0_en];
      Register_inst187 <= _T_190[_T_2 == 8'hBB & write_0_en];
      Register_inst188 <= _T_191[_T_2 == 8'hBC & write_0_en];
      Register_inst189 <= _T_192[_T_2 == 8'hBD & write_0_en];
      Register_inst190 <= _T_193[_T_2 == 8'hBE & write_0_en];
      Register_inst191 <= _T_194[_T_2 == 8'hBF & write_0_en];
      Register_inst192 <= _T_195[_T_2 == 8'hC0 & write_0_en];
      Register_inst193 <= _T_196[_T_2 == 8'hC1 & write_0_en];
      Register_inst194 <= _T_197[_T_2 == 8'hC2 & write_0_en];
      Register_inst195 <= _T_198[_T_2 == 8'hC3 & write_0_en];
      Register_inst196 <= _T_199[_T_2 == 8'hC4 & write_0_en];
      Register_inst197 <= _T_200[_T_2 == 8'hC5 & write_0_en];
      Register_inst198 <= _T_201[_T_2 == 8'hC6 & write_0_en];
      Register_inst199 <= _T_202[_T_2 == 8'hC7 & write_0_en];
      Register_inst200 <= _T_203[_T_2 == 8'hC8 & write_0_en];
      Register_inst201 <= _T_204[_T_2 == 8'hC9 & write_0_en];
      Register_inst202 <= _T_205[_T_2 == 8'hCA & write_0_en];
      Register_inst203 <= _T_206[_T_2 == 8'hCB & write_0_en];
      Register_inst204 <= _T_207[_T_2 == 8'hCC & write_0_en];
      Register_inst205 <= _T_208[_T_2 == 8'hCD & write_0_en];
      Register_inst206 <= _T_209[_T_2 == 8'hCE & write_0_en];
      Register_inst207 <= _T_210[_T_2 == 8'hCF & write_0_en];
      Register_inst208 <= _T_211[_T_2 == 8'hD0 & write_0_en];
      Register_inst209 <= _T_212[_T_2 == 8'hD1 & write_0_en];
      Register_inst210 <= _T_213[_T_2 == 8'hD2 & write_0_en];
      Register_inst211 <= _T_214[_T_2 == 8'hD3 & write_0_en];
      Register_inst212 <= _T_215[_T_2 == 8'hD4 & write_0_en];
      Register_inst213 <= _T_216[_T_2 == 8'hD5 & write_0_en];
      Register_inst214 <= _T_217[_T_2 == 8'hD6 & write_0_en];
      Register_inst215 <= _T_218[_T_2 == 8'hD7 & write_0_en];
      Register_inst216 <= _T_219[_T_2 == 8'hD8 & write_0_en];
      Register_inst217 <= _T_220[_T_2 == 8'hD9 & write_0_en];
      Register_inst218 <= _T_221[_T_2 == 8'hDA & write_0_en];
      Register_inst219 <= _T_222[_T_2 == 8'hDB & write_0_en];
      Register_inst220 <= _T_223[_T_2 == 8'hDC & write_0_en];
      Register_inst221 <= _T_224[_T_2 == 8'hDD & write_0_en];
      Register_inst222 <= _T_225[_T_2 == 8'hDE & write_0_en];
      Register_inst223 <= _T_226[_T_2 == 8'hDF & write_0_en];
      Register_inst224 <= _T_227[_T_2 == 8'hE0 & write_0_en];
      Register_inst225 <= _T_228[_T_2 == 8'hE1 & write_0_en];
      Register_inst226 <= _T_229[_T_2 == 8'hE2 & write_0_en];
      Register_inst227 <= _T_230[_T_2 == 8'hE3 & write_0_en];
      Register_inst228 <= _T_231[_T_2 == 8'hE4 & write_0_en];
      Register_inst229 <= _T_232[_T_2 == 8'hE5 & write_0_en];
      Register_inst230 <= _T_233[_T_2 == 8'hE6 & write_0_en];
      Register_inst231 <= _T_234[_T_2 == 8'hE7 & write_0_en];
      Register_inst232 <= _T_235[_T_2 == 8'hE8 & write_0_en];
      Register_inst233 <= _T_236[_T_2 == 8'hE9 & write_0_en];
      Register_inst234 <= _T_237[_T_2 == 8'hEA & write_0_en];
      Register_inst235 <= _T_238[_T_2 == 8'hEB & write_0_en];
      Register_inst236 <= _T_239[_T_2 == 8'hEC & write_0_en];
      Register_inst237 <= _T_240[_T_2 == 8'hED & write_0_en];
      Register_inst238 <= _T_241[_T_2 == 8'hEE & write_0_en];
      Register_inst239 <= _T_242[_T_2 == 8'hEF & write_0_en];
      Register_inst240 <= _T_243[_T_2 == 8'hF0 & write_0_en];
      Register_inst241 <= _T_244[_T_2 == 8'hF1 & write_0_en];
      Register_inst242 <= _T_245[_T_2 == 8'hF2 & write_0_en];
      Register_inst243 <= _T_246[_T_2 == 8'hF3 & write_0_en];
      Register_inst244 <= _T_247[_T_2 == 8'hF4 & write_0_en];
      Register_inst245 <= _T_248[_T_2 == 8'hF5 & write_0_en];
      Register_inst246 <= _T_249[_T_2 == 8'hF6 & write_0_en];
      Register_inst247 <= _T_250[_T_2 == 8'hF7 & write_0_en];
      Register_inst248 <= _T_251[_T_2 == 8'hF8 & write_0_en];
      Register_inst249 <= _T_252[_T_2 == 8'hF9 & write_0_en];
      Register_inst250 <= _T_253[_T_2 == 8'hFA & write_0_en];
      Register_inst251 <= _T_254[_T_2 == 8'hFB & write_0_en];
      Register_inst252 <= _T_255[_T_2 == 8'hFC & write_0_en];
      Register_inst253 <= _T_256[_T_2 == 8'hFD & write_0_en];
      Register_inst254 <= _T_257[_T_2 == 8'hFE & write_0_en];
      Register_inst255 <= _T_258[&_T_2 & write_0_en];
    end
  end // always_ff @(posedge or posedge)
  initial begin
    Register_inst0 = 32'h0;
    Register_inst1 = 32'h0;
    Register_inst2 = 32'h0;
    Register_inst3 = 32'h0;
    Register_inst4 = 32'h0;
    Register_inst5 = 32'h0;
    Register_inst6 = 32'h0;
    Register_inst7 = 32'h0;
    Register_inst8 = 32'h0;
    Register_inst9 = 32'h0;
    Register_inst10 = 32'h0;
    Register_inst11 = 32'h0;
    Register_inst12 = 32'h0;
    Register_inst13 = 32'h0;
    Register_inst14 = 32'h0;
    Register_inst15 = 32'h0;
    Register_inst16 = 32'h0;
    Register_inst17 = 32'h0;
    Register_inst18 = 32'h0;
    Register_inst19 = 32'h0;
    Register_inst20 = 32'h0;
    Register_inst21 = 32'h0;
    Register_inst22 = 32'h0;
    Register_inst23 = 32'h0;
    Register_inst24 = 32'h0;
    Register_inst25 = 32'h0;
    Register_inst26 = 32'h0;
    Register_inst27 = 32'h0;
    Register_inst28 = 32'h0;
    Register_inst29 = 32'h0;
    Register_inst30 = 32'h0;
    Register_inst31 = 32'h0;
    Register_inst32 = 32'h0;
    Register_inst33 = 32'h0;
    Register_inst34 = 32'h0;
    Register_inst35 = 32'h0;
    Register_inst36 = 32'h0;
    Register_inst37 = 32'h0;
    Register_inst38 = 32'h0;
    Register_inst39 = 32'h0;
    Register_inst40 = 32'h0;
    Register_inst41 = 32'h0;
    Register_inst42 = 32'h0;
    Register_inst43 = 32'h0;
    Register_inst44 = 32'h0;
    Register_inst45 = 32'h0;
    Register_inst46 = 32'h0;
    Register_inst47 = 32'h0;
    Register_inst48 = 32'h0;
    Register_inst49 = 32'h0;
    Register_inst50 = 32'h0;
    Register_inst51 = 32'h0;
    Register_inst52 = 32'h0;
    Register_inst53 = 32'h0;
    Register_inst54 = 32'h0;
    Register_inst55 = 32'h0;
    Register_inst56 = 32'h0;
    Register_inst57 = 32'h0;
    Register_inst58 = 32'h0;
    Register_inst59 = 32'h0;
    Register_inst60 = 32'h0;
    Register_inst61 = 32'h0;
    Register_inst62 = 32'h0;
    Register_inst63 = 32'h0;
    Register_inst64 = 32'h0;
    Register_inst65 = 32'h0;
    Register_inst66 = 32'h0;
    Register_inst67 = 32'h0;
    Register_inst68 = 32'h0;
    Register_inst69 = 32'h0;
    Register_inst70 = 32'h0;
    Register_inst71 = 32'h0;
    Register_inst72 = 32'h0;
    Register_inst73 = 32'h0;
    Register_inst74 = 32'h0;
    Register_inst75 = 32'h0;
    Register_inst76 = 32'h0;
    Register_inst77 = 32'h0;
    Register_inst78 = 32'h0;
    Register_inst79 = 32'h0;
    Register_inst80 = 32'h0;
    Register_inst81 = 32'h0;
    Register_inst82 = 32'h0;
    Register_inst83 = 32'h0;
    Register_inst84 = 32'h0;
    Register_inst85 = 32'h0;
    Register_inst86 = 32'h0;
    Register_inst87 = 32'h0;
    Register_inst88 = 32'h0;
    Register_inst89 = 32'h0;
    Register_inst90 = 32'h0;
    Register_inst91 = 32'h0;
    Register_inst92 = 32'h0;
    Register_inst93 = 32'h0;
    Register_inst94 = 32'h0;
    Register_inst95 = 32'h0;
    Register_inst96 = 32'h0;
    Register_inst97 = 32'h0;
    Register_inst98 = 32'h0;
    Register_inst99 = 32'h0;
    Register_inst100 = 32'h0;
    Register_inst101 = 32'h0;
    Register_inst102 = 32'h0;
    Register_inst103 = 32'h0;
    Register_inst104 = 32'h0;
    Register_inst105 = 32'h0;
    Register_inst106 = 32'h0;
    Register_inst107 = 32'h0;
    Register_inst108 = 32'h0;
    Register_inst109 = 32'h0;
    Register_inst110 = 32'h0;
    Register_inst111 = 32'h0;
    Register_inst112 = 32'h0;
    Register_inst113 = 32'h0;
    Register_inst114 = 32'h0;
    Register_inst115 = 32'h0;
    Register_inst116 = 32'h0;
    Register_inst117 = 32'h0;
    Register_inst118 = 32'h0;
    Register_inst119 = 32'h0;
    Register_inst120 = 32'h0;
    Register_inst121 = 32'h0;
    Register_inst122 = 32'h0;
    Register_inst123 = 32'h0;
    Register_inst124 = 32'h0;
    Register_inst125 = 32'h0;
    Register_inst126 = 32'h0;
    Register_inst127 = 32'h0;
    Register_inst128 = 32'h0;
    Register_inst129 = 32'h0;
    Register_inst130 = 32'h0;
    Register_inst131 = 32'h0;
    Register_inst132 = 32'h0;
    Register_inst133 = 32'h0;
    Register_inst134 = 32'h0;
    Register_inst135 = 32'h0;
    Register_inst136 = 32'h0;
    Register_inst137 = 32'h0;
    Register_inst138 = 32'h0;
    Register_inst139 = 32'h0;
    Register_inst140 = 32'h0;
    Register_inst141 = 32'h0;
    Register_inst142 = 32'h0;
    Register_inst143 = 32'h0;
    Register_inst144 = 32'h0;
    Register_inst145 = 32'h0;
    Register_inst146 = 32'h0;
    Register_inst147 = 32'h0;
    Register_inst148 = 32'h0;
    Register_inst149 = 32'h0;
    Register_inst150 = 32'h0;
    Register_inst151 = 32'h0;
    Register_inst152 = 32'h0;
    Register_inst153 = 32'h0;
    Register_inst154 = 32'h0;
    Register_inst155 = 32'h0;
    Register_inst156 = 32'h0;
    Register_inst157 = 32'h0;
    Register_inst158 = 32'h0;
    Register_inst159 = 32'h0;
    Register_inst160 = 32'h0;
    Register_inst161 = 32'h0;
    Register_inst162 = 32'h0;
    Register_inst163 = 32'h0;
    Register_inst164 = 32'h0;
    Register_inst165 = 32'h0;
    Register_inst166 = 32'h0;
    Register_inst167 = 32'h0;
    Register_inst168 = 32'h0;
    Register_inst169 = 32'h0;
    Register_inst170 = 32'h0;
    Register_inst171 = 32'h0;
    Register_inst172 = 32'h0;
    Register_inst173 = 32'h0;
    Register_inst174 = 32'h0;
    Register_inst175 = 32'h0;
    Register_inst176 = 32'h0;
    Register_inst177 = 32'h0;
    Register_inst178 = 32'h0;
    Register_inst179 = 32'h0;
    Register_inst180 = 32'h0;
    Register_inst181 = 32'h0;
    Register_inst182 = 32'h0;
    Register_inst183 = 32'h0;
    Register_inst184 = 32'h0;
    Register_inst185 = 32'h0;
    Register_inst186 = 32'h0;
    Register_inst187 = 32'h0;
    Register_inst188 = 32'h0;
    Register_inst189 = 32'h0;
    Register_inst190 = 32'h0;
    Register_inst191 = 32'h0;
    Register_inst192 = 32'h0;
    Register_inst193 = 32'h0;
    Register_inst194 = 32'h0;
    Register_inst195 = 32'h0;
    Register_inst196 = 32'h0;
    Register_inst197 = 32'h0;
    Register_inst198 = 32'h0;
    Register_inst199 = 32'h0;
    Register_inst200 = 32'h0;
    Register_inst201 = 32'h0;
    Register_inst202 = 32'h0;
    Register_inst203 = 32'h0;
    Register_inst204 = 32'h0;
    Register_inst205 = 32'h0;
    Register_inst206 = 32'h0;
    Register_inst207 = 32'h0;
    Register_inst208 = 32'h0;
    Register_inst209 = 32'h0;
    Register_inst210 = 32'h0;
    Register_inst211 = 32'h0;
    Register_inst212 = 32'h0;
    Register_inst213 = 32'h0;
    Register_inst214 = 32'h0;
    Register_inst215 = 32'h0;
    Register_inst216 = 32'h0;
    Register_inst217 = 32'h0;
    Register_inst218 = 32'h0;
    Register_inst219 = 32'h0;
    Register_inst220 = 32'h0;
    Register_inst221 = 32'h0;
    Register_inst222 = 32'h0;
    Register_inst223 = 32'h0;
    Register_inst224 = 32'h0;
    Register_inst225 = 32'h0;
    Register_inst226 = 32'h0;
    Register_inst227 = 32'h0;
    Register_inst228 = 32'h0;
    Register_inst229 = 32'h0;
    Register_inst230 = 32'h0;
    Register_inst231 = 32'h0;
    Register_inst232 = 32'h0;
    Register_inst233 = 32'h0;
    Register_inst234 = 32'h0;
    Register_inst235 = 32'h0;
    Register_inst236 = 32'h0;
    Register_inst237 = 32'h0;
    Register_inst238 = 32'h0;
    Register_inst239 = 32'h0;
    Register_inst240 = 32'h0;
    Register_inst241 = 32'h0;
    Register_inst242 = 32'h0;
    Register_inst243 = 32'h0;
    Register_inst244 = 32'h0;
    Register_inst245 = 32'h0;
    Register_inst246 = 32'h0;
    Register_inst247 = 32'h0;
    Register_inst248 = 32'h0;
    Register_inst249 = 32'h0;
    Register_inst250 = 32'h0;
    Register_inst251 = 32'h0;
    Register_inst252 = 32'h0;
    Register_inst253 = 32'h0;
    Register_inst254 = 32'h0;
    Register_inst255 = 32'h0;
  end // initial
  wire [255:0][31:0] _T = {{Register_inst0}, {Register_inst1}, {Register_inst2}, {Register_inst3}, {Register_inst4},
                {Register_inst5}, {Register_inst6}, {Register_inst7}, {Register_inst8}, {Register_inst9},
                {Register_inst10}, {Register_inst11}, {Register_inst12}, {Register_inst13},
                {Register_inst14}, {Register_inst15}, {Register_inst16}, {Register_inst17},
                {Register_inst18}, {Register_inst19}, {Register_inst20}, {Register_inst21},
                {Register_inst22}, {Register_inst23}, {Register_inst24}, {Register_inst25},
                {Register_inst26}, {Register_inst27}, {Register_inst28}, {Register_inst29},
                {Register_inst30}, {Register_inst31}, {Register_inst32}, {Register_inst33},
                {Register_inst34}, {Register_inst35}, {Register_inst36}, {Register_inst37},
                {Register_inst38}, {Register_inst39}, {Register_inst40}, {Register_inst41},
                {Register_inst42}, {Register_inst43}, {Register_inst44}, {Register_inst45},
                {Register_inst46}, {Register_inst47}, {Register_inst48}, {Register_inst49},
                {Register_inst50}, {Register_inst51}, {Register_inst52}, {Register_inst53},
                {Register_inst54}, {Register_inst55}, {Register_inst56}, {Register_inst57},
                {Register_inst58}, {Register_inst59}, {Register_inst60}, {Register_inst61},
                {Register_inst62}, {Register_inst63}, {Register_inst64}, {Register_inst65},
                {Register_inst66}, {Register_inst67}, {Register_inst68}, {Register_inst69},
                {Register_inst70}, {Register_inst71}, {Register_inst72}, {Register_inst73},
                {Register_inst74}, {Register_inst75}, {Register_inst76}, {Register_inst77},
                {Register_inst78}, {Register_inst79}, {Register_inst80}, {Register_inst81},
                {Register_inst82}, {Register_inst83}, {Register_inst84}, {Register_inst85},
                {Register_inst86}, {Register_inst87}, {Register_inst88}, {Register_inst89},
                {Register_inst90}, {Register_inst91}, {Register_inst92}, {Register_inst93},
                {Register_inst94}, {Register_inst95}, {Register_inst96}, {Register_inst97},
                {Register_inst98}, {Register_inst99}, {Register_inst100}, {Register_inst101},
                {Register_inst102}, {Register_inst103}, {Register_inst104}, {Register_inst105},
                {Register_inst106}, {Register_inst107}, {Register_inst108}, {Register_inst109},
                {Register_inst110}, {Register_inst111}, {Register_inst112}, {Register_inst113},
                {Register_inst114}, {Register_inst115}, {Register_inst116}, {Register_inst117},
                {Register_inst118}, {Register_inst119}, {Register_inst120}, {Register_inst121},
                {Register_inst122}, {Register_inst123}, {Register_inst124}, {Register_inst125},
                {Register_inst126}, {Register_inst127}, {Register_inst128}, {Register_inst129},
                {Register_inst130}, {Register_inst131}, {Register_inst132}, {Register_inst133},
                {Register_inst134}, {Register_inst135}, {Register_inst136}, {Register_inst137},
                {Register_inst138}, {Register_inst139}, {Register_inst140}, {Register_inst141},
                {Register_inst142}, {Register_inst143}, {Register_inst144}, {Register_inst145},
                {Register_inst146}, {Register_inst147}, {Register_inst148}, {Register_inst149},
                {Register_inst150}, {Register_inst151}, {Register_inst152}, {Register_inst153},
                {Register_inst154}, {Register_inst155}, {Register_inst156}, {Register_inst157},
                {Register_inst158}, {Register_inst159}, {Register_inst160}, {Register_inst161},
                {Register_inst162}, {Register_inst163}, {Register_inst164}, {Register_inst165},
                {Register_inst166}, {Register_inst167}, {Register_inst168}, {Register_inst169},
                {Register_inst170}, {Register_inst171}, {Register_inst172}, {Register_inst173},
                {Register_inst174}, {Register_inst175}, {Register_inst176}, {Register_inst177},
                {Register_inst178}, {Register_inst179}, {Register_inst180}, {Register_inst181},
                {Register_inst182}, {Register_inst183}, {Register_inst184}, {Register_inst185},
                {Register_inst186}, {Register_inst187}, {Register_inst188}, {Register_inst189},
                {Register_inst190}, {Register_inst191}, {Register_inst192}, {Register_inst193},
                {Register_inst194}, {Register_inst195}, {Register_inst196}, {Register_inst197},
                {Register_inst198}, {Register_inst199}, {Register_inst200}, {Register_inst201},
                {Register_inst202}, {Register_inst203}, {Register_inst204}, {Register_inst205},
                {Register_inst206}, {Register_inst207}, {Register_inst208}, {Register_inst209},
                {Register_inst210}, {Register_inst211}, {Register_inst212}, {Register_inst213},
                {Register_inst214}, {Register_inst215}, {Register_inst216}, {Register_inst217},
                {Register_inst218}, {Register_inst219}, {Register_inst220}, {Register_inst221},
                {Register_inst222}, {Register_inst223}, {Register_inst224}, {Register_inst225},
                {Register_inst226}, {Register_inst227}, {Register_inst228}, {Register_inst229},
                {Register_inst230}, {Register_inst231}, {Register_inst232}, {Register_inst233},
                {Register_inst234}, {Register_inst235}, {Register_inst236}, {Register_inst237},
                {Register_inst238}, {Register_inst239}, {Register_inst240}, {Register_inst241},
                {Register_inst242}, {Register_inst243}, {Register_inst244}, {Register_inst245},
                {Register_inst246}, {Register_inst247}, {Register_inst248}, {Register_inst249},
                {Register_inst250}, {Register_inst251}, {Register_inst252}, {Register_inst253},
                {Register_inst254}, {Register_inst255}};
  wire [255:0][31:0] _T_0 = {{Register_inst0}, {Register_inst1}, {Register_inst2}, {Register_inst3}, {Register_inst4},
                {Register_inst5}, {Register_inst6}, {Register_inst7}, {Register_inst8}, {Register_inst9},
                {Register_inst10}, {Register_inst11}, {Register_inst12}, {Register_inst13},
                {Register_inst14}, {Register_inst15}, {Register_inst16}, {Register_inst17},
                {Register_inst18}, {Register_inst19}, {Register_inst20}, {Register_inst21},
                {Register_inst22}, {Register_inst23}, {Register_inst24}, {Register_inst25},
                {Register_inst26}, {Register_inst27}, {Register_inst28}, {Register_inst29},
                {Register_inst30}, {Register_inst31}, {Register_inst32}, {Register_inst33},
                {Register_inst34}, {Register_inst35}, {Register_inst36}, {Register_inst37},
                {Register_inst38}, {Register_inst39}, {Register_inst40}, {Register_inst41},
                {Register_inst42}, {Register_inst43}, {Register_inst44}, {Register_inst45},
                {Register_inst46}, {Register_inst47}, {Register_inst48}, {Register_inst49},
                {Register_inst50}, {Register_inst51}, {Register_inst52}, {Register_inst53},
                {Register_inst54}, {Register_inst55}, {Register_inst56}, {Register_inst57},
                {Register_inst58}, {Register_inst59}, {Register_inst60}, {Register_inst61},
                {Register_inst62}, {Register_inst63}, {Register_inst64}, {Register_inst65},
                {Register_inst66}, {Register_inst67}, {Register_inst68}, {Register_inst69},
                {Register_inst70}, {Register_inst71}, {Register_inst72}, {Register_inst73},
                {Register_inst74}, {Register_inst75}, {Register_inst76}, {Register_inst77},
                {Register_inst78}, {Register_inst79}, {Register_inst80}, {Register_inst81},
                {Register_inst82}, {Register_inst83}, {Register_inst84}, {Register_inst85},
                {Register_inst86}, {Register_inst87}, {Register_inst88}, {Register_inst89},
                {Register_inst90}, {Register_inst91}, {Register_inst92}, {Register_inst93},
                {Register_inst94}, {Register_inst95}, {Register_inst96}, {Register_inst97},
                {Register_inst98}, {Register_inst99}, {Register_inst100}, {Register_inst101},
                {Register_inst102}, {Register_inst103}, {Register_inst104}, {Register_inst105},
                {Register_inst106}, {Register_inst107}, {Register_inst108}, {Register_inst109},
                {Register_inst110}, {Register_inst111}, {Register_inst112}, {Register_inst113},
                {Register_inst114}, {Register_inst115}, {Register_inst116}, {Register_inst117},
                {Register_inst118}, {Register_inst119}, {Register_inst120}, {Register_inst121},
                {Register_inst122}, {Register_inst123}, {Register_inst124}, {Register_inst125},
                {Register_inst126}, {Register_inst127}, {Register_inst128}, {Register_inst129},
                {Register_inst130}, {Register_inst131}, {Register_inst132}, {Register_inst133},
                {Register_inst134}, {Register_inst135}, {Register_inst136}, {Register_inst137},
                {Register_inst138}, {Register_inst139}, {Register_inst140}, {Register_inst141},
                {Register_inst142}, {Register_inst143}, {Register_inst144}, {Register_inst145},
                {Register_inst146}, {Register_inst147}, {Register_inst148}, {Register_inst149},
                {Register_inst150}, {Register_inst151}, {Register_inst152}, {Register_inst153},
                {Register_inst154}, {Register_inst155}, {Register_inst156}, {Register_inst157},
                {Register_inst158}, {Register_inst159}, {Register_inst160}, {Register_inst161},
                {Register_inst162}, {Register_inst163}, {Register_inst164}, {Register_inst165},
                {Register_inst166}, {Register_inst167}, {Register_inst168}, {Register_inst169},
                {Register_inst170}, {Register_inst171}, {Register_inst172}, {Register_inst173},
                {Register_inst174}, {Register_inst175}, {Register_inst176}, {Register_inst177},
                {Register_inst178}, {Register_inst179}, {Register_inst180}, {Register_inst181},
                {Register_inst182}, {Register_inst183}, {Register_inst184}, {Register_inst185},
                {Register_inst186}, {Register_inst187}, {Register_inst188}, {Register_inst189},
                {Register_inst190}, {Register_inst191}, {Register_inst192}, {Register_inst193},
                {Register_inst194}, {Register_inst195}, {Register_inst196}, {Register_inst197},
                {Register_inst198}, {Register_inst199}, {Register_inst200}, {Register_inst201},
                {Register_inst202}, {Register_inst203}, {Register_inst204}, {Register_inst205},
                {Register_inst206}, {Register_inst207}, {Register_inst208}, {Register_inst209},
                {Register_inst210}, {Register_inst211}, {Register_inst212}, {Register_inst213},
                {Register_inst214}, {Register_inst215}, {Register_inst216}, {Register_inst217},
                {Register_inst218}, {Register_inst219}, {Register_inst220}, {Register_inst221},
                {Register_inst222}, {Register_inst223}, {Register_inst224}, {Register_inst225},
                {Register_inst226}, {Register_inst227}, {Register_inst228}, {Register_inst229},
                {Register_inst230}, {Register_inst231}, {Register_inst232}, {Register_inst233},
                {Register_inst234}, {Register_inst235}, {Register_inst236}, {Register_inst237},
                {Register_inst238}, {Register_inst239}, {Register_inst240}, {Register_inst241},
                {Register_inst242}, {Register_inst243}, {Register_inst244}, {Register_inst245},
                {Register_inst246}, {Register_inst247}, {Register_inst248}, {Register_inst249},
                {Register_inst250}, {Register_inst251}, {Register_inst252}, {Register_inst253},
                {Register_inst254}, {Register_inst255}};
  assign file_read_0_data = _T[file_read_0_addr];
  assign file_read_1_data = _T_0[file_read_1_addr];
endmodule

module code(
  input                                                        CLK, ASYNCRESET,
  input  [7:0]                                                 code_read_0_addr,
  input  struct packed {logic [31:0] data; logic [7:0] addr; } write_0,
  input                                                        write_0_en,
  output [31:0]                                                code_read_0_data);

  reg [31:0] Register_inst0;
  reg [31:0] Register_inst1;
  reg [31:0] Register_inst2;
  reg [31:0] Register_inst3;
  reg [31:0] Register_inst4;
  reg [31:0] Register_inst5;
  reg [31:0] Register_inst6;
  reg [31:0] Register_inst7;
  reg [31:0] Register_inst8;
  reg [31:0] Register_inst9;
  reg [31:0] Register_inst10;
  reg [31:0] Register_inst11;
  reg [31:0] Register_inst12;
  reg [31:0] Register_inst13;
  reg [31:0] Register_inst14;
  reg [31:0] Register_inst15;
  reg [31:0] Register_inst16;
  reg [31:0] Register_inst17;
  reg [31:0] Register_inst18;
  reg [31:0] Register_inst19;
  reg [31:0] Register_inst20;
  reg [31:0] Register_inst21;
  reg [31:0] Register_inst22;
  reg [31:0] Register_inst23;
  reg [31:0] Register_inst24;
  reg [31:0] Register_inst25;
  reg [31:0] Register_inst26;
  reg [31:0] Register_inst27;
  reg [31:0] Register_inst28;
  reg [31:0] Register_inst29;
  reg [31:0] Register_inst30;
  reg [31:0] Register_inst31;
  reg [31:0] Register_inst32;
  reg [31:0] Register_inst33;
  reg [31:0] Register_inst34;
  reg [31:0] Register_inst35;
  reg [31:0] Register_inst36;
  reg [31:0] Register_inst37;
  reg [31:0] Register_inst38;
  reg [31:0] Register_inst39;
  reg [31:0] Register_inst40;
  reg [31:0] Register_inst41;
  reg [31:0] Register_inst42;
  reg [31:0] Register_inst43;
  reg [31:0] Register_inst44;
  reg [31:0] Register_inst45;
  reg [31:0] Register_inst46;
  reg [31:0] Register_inst47;
  reg [31:0] Register_inst48;
  reg [31:0] Register_inst49;
  reg [31:0] Register_inst50;
  reg [31:0] Register_inst51;
  reg [31:0] Register_inst52;
  reg [31:0] Register_inst53;
  reg [31:0] Register_inst54;
  reg [31:0] Register_inst55;
  reg [31:0] Register_inst56;
  reg [31:0] Register_inst57;
  reg [31:0] Register_inst58;
  reg [31:0] Register_inst59;
  reg [31:0] Register_inst60;
  reg [31:0] Register_inst61;
  reg [31:0] Register_inst62;
  reg [31:0] Register_inst63;
  reg [31:0] Register_inst64;
  reg [31:0] Register_inst65;
  reg [31:0] Register_inst66;
  reg [31:0] Register_inst67;
  reg [31:0] Register_inst68;
  reg [31:0] Register_inst69;
  reg [31:0] Register_inst70;
  reg [31:0] Register_inst71;
  reg [31:0] Register_inst72;
  reg [31:0] Register_inst73;
  reg [31:0] Register_inst74;
  reg [31:0] Register_inst75;
  reg [31:0] Register_inst76;
  reg [31:0] Register_inst77;
  reg [31:0] Register_inst78;
  reg [31:0] Register_inst79;
  reg [31:0] Register_inst80;
  reg [31:0] Register_inst81;
  reg [31:0] Register_inst82;
  reg [31:0] Register_inst83;
  reg [31:0] Register_inst84;
  reg [31:0] Register_inst85;
  reg [31:0] Register_inst86;
  reg [31:0] Register_inst87;
  reg [31:0] Register_inst88;
  reg [31:0] Register_inst89;
  reg [31:0] Register_inst90;
  reg [31:0] Register_inst91;
  reg [31:0] Register_inst92;
  reg [31:0] Register_inst93;
  reg [31:0] Register_inst94;
  reg [31:0] Register_inst95;
  reg [31:0] Register_inst96;
  reg [31:0] Register_inst97;
  reg [31:0] Register_inst98;
  reg [31:0] Register_inst99;
  reg [31:0] Register_inst100;
  reg [31:0] Register_inst101;
  reg [31:0] Register_inst102;
  reg [31:0] Register_inst103;
  reg [31:0] Register_inst104;
  reg [31:0] Register_inst105;
  reg [31:0] Register_inst106;
  reg [31:0] Register_inst107;
  reg [31:0] Register_inst108;
  reg [31:0] Register_inst109;
  reg [31:0] Register_inst110;
  reg [31:0] Register_inst111;
  reg [31:0] Register_inst112;
  reg [31:0] Register_inst113;
  reg [31:0] Register_inst114;
  reg [31:0] Register_inst115;
  reg [31:0] Register_inst116;
  reg [31:0] Register_inst117;
  reg [31:0] Register_inst118;
  reg [31:0] Register_inst119;
  reg [31:0] Register_inst120;
  reg [31:0] Register_inst121;
  reg [31:0] Register_inst122;
  reg [31:0] Register_inst123;
  reg [31:0] Register_inst124;
  reg [31:0] Register_inst125;
  reg [31:0] Register_inst126;
  reg [31:0] Register_inst127;
  reg [31:0] Register_inst128;
  reg [31:0] Register_inst129;
  reg [31:0] Register_inst130;
  reg [31:0] Register_inst131;
  reg [31:0] Register_inst132;
  reg [31:0] Register_inst133;
  reg [31:0] Register_inst134;
  reg [31:0] Register_inst135;
  reg [31:0] Register_inst136;
  reg [31:0] Register_inst137;
  reg [31:0] Register_inst138;
  reg [31:0] Register_inst139;
  reg [31:0] Register_inst140;
  reg [31:0] Register_inst141;
  reg [31:0] Register_inst142;
  reg [31:0] Register_inst143;
  reg [31:0] Register_inst144;
  reg [31:0] Register_inst145;
  reg [31:0] Register_inst146;
  reg [31:0] Register_inst147;
  reg [31:0] Register_inst148;
  reg [31:0] Register_inst149;
  reg [31:0] Register_inst150;
  reg [31:0] Register_inst151;
  reg [31:0] Register_inst152;
  reg [31:0] Register_inst153;
  reg [31:0] Register_inst154;
  reg [31:0] Register_inst155;
  reg [31:0] Register_inst156;
  reg [31:0] Register_inst157;
  reg [31:0] Register_inst158;
  reg [31:0] Register_inst159;
  reg [31:0] Register_inst160;
  reg [31:0] Register_inst161;
  reg [31:0] Register_inst162;
  reg [31:0] Register_inst163;
  reg [31:0] Register_inst164;
  reg [31:0] Register_inst165;
  reg [31:0] Register_inst166;
  reg [31:0] Register_inst167;
  reg [31:0] Register_inst168;
  reg [31:0] Register_inst169;
  reg [31:0] Register_inst170;
  reg [31:0] Register_inst171;
  reg [31:0] Register_inst172;
  reg [31:0] Register_inst173;
  reg [31:0] Register_inst174;
  reg [31:0] Register_inst175;
  reg [31:0] Register_inst176;
  reg [31:0] Register_inst177;
  reg [31:0] Register_inst178;
  reg [31:0] Register_inst179;
  reg [31:0] Register_inst180;
  reg [31:0] Register_inst181;
  reg [31:0] Register_inst182;
  reg [31:0] Register_inst183;
  reg [31:0] Register_inst184;
  reg [31:0] Register_inst185;
  reg [31:0] Register_inst186;
  reg [31:0] Register_inst187;
  reg [31:0] Register_inst188;
  reg [31:0] Register_inst189;
  reg [31:0] Register_inst190;
  reg [31:0] Register_inst191;
  reg [31:0] Register_inst192;
  reg [31:0] Register_inst193;
  reg [31:0] Register_inst194;
  reg [31:0] Register_inst195;
  reg [31:0] Register_inst196;
  reg [31:0] Register_inst197;
  reg [31:0] Register_inst198;
  reg [31:0] Register_inst199;
  reg [31:0] Register_inst200;
  reg [31:0] Register_inst201;
  reg [31:0] Register_inst202;
  reg [31:0] Register_inst203;
  reg [31:0] Register_inst204;
  reg [31:0] Register_inst205;
  reg [31:0] Register_inst206;
  reg [31:0] Register_inst207;
  reg [31:0] Register_inst208;
  reg [31:0] Register_inst209;
  reg [31:0] Register_inst210;
  reg [31:0] Register_inst211;
  reg [31:0] Register_inst212;
  reg [31:0] Register_inst213;
  reg [31:0] Register_inst214;
  reg [31:0] Register_inst215;
  reg [31:0] Register_inst216;
  reg [31:0] Register_inst217;
  reg [31:0] Register_inst218;
  reg [31:0] Register_inst219;
  reg [31:0] Register_inst220;
  reg [31:0] Register_inst221;
  reg [31:0] Register_inst222;
  reg [31:0] Register_inst223;
  reg [31:0] Register_inst224;
  reg [31:0] Register_inst225;
  reg [31:0] Register_inst226;
  reg [31:0] Register_inst227;
  reg [31:0] Register_inst228;
  reg [31:0] Register_inst229;
  reg [31:0] Register_inst230;
  reg [31:0] Register_inst231;
  reg [31:0] Register_inst232;
  reg [31:0] Register_inst233;
  reg [31:0] Register_inst234;
  reg [31:0] Register_inst235;
  reg [31:0] Register_inst236;
  reg [31:0] Register_inst237;
  reg [31:0] Register_inst238;
  reg [31:0] Register_inst239;
  reg [31:0] Register_inst240;
  reg [31:0] Register_inst241;
  reg [31:0] Register_inst242;
  reg [31:0] Register_inst243;
  reg [31:0] Register_inst244;
  reg [31:0] Register_inst245;
  reg [31:0] Register_inst246;
  reg [31:0] Register_inst247;
  reg [31:0] Register_inst248;
  reg [31:0] Register_inst249;
  reg [31:0] Register_inst250;
  reg [31:0] Register_inst251;
  reg [31:0] Register_inst252;
  reg [31:0] Register_inst253;
  reg [31:0] Register_inst254;
  reg [31:0] Register_inst255;

  always_ff @(posedge CLK or posedge ASYNCRESET) begin
    if (ASYNCRESET) begin
      Register_inst0 <= 32'h0;
      Register_inst1 <= 32'h0;
      Register_inst2 <= 32'h0;
      Register_inst3 <= 32'h0;
      Register_inst4 <= 32'h0;
      Register_inst5 <= 32'h0;
      Register_inst6 <= 32'h0;
      Register_inst7 <= 32'h0;
      Register_inst8 <= 32'h0;
      Register_inst9 <= 32'h0;
      Register_inst10 <= 32'h0;
      Register_inst11 <= 32'h0;
      Register_inst12 <= 32'h0;
      Register_inst13 <= 32'h0;
      Register_inst14 <= 32'h0;
      Register_inst15 <= 32'h0;
      Register_inst16 <= 32'h0;
      Register_inst17 <= 32'h0;
      Register_inst18 <= 32'h0;
      Register_inst19 <= 32'h0;
      Register_inst20 <= 32'h0;
      Register_inst21 <= 32'h0;
      Register_inst22 <= 32'h0;
      Register_inst23 <= 32'h0;
      Register_inst24 <= 32'h0;
      Register_inst25 <= 32'h0;
      Register_inst26 <= 32'h0;
      Register_inst27 <= 32'h0;
      Register_inst28 <= 32'h0;
      Register_inst29 <= 32'h0;
      Register_inst30 <= 32'h0;
      Register_inst31 <= 32'h0;
      Register_inst32 <= 32'h0;
      Register_inst33 <= 32'h0;
      Register_inst34 <= 32'h0;
      Register_inst35 <= 32'h0;
      Register_inst36 <= 32'h0;
      Register_inst37 <= 32'h0;
      Register_inst38 <= 32'h0;
      Register_inst39 <= 32'h0;
      Register_inst40 <= 32'h0;
      Register_inst41 <= 32'h0;
      Register_inst42 <= 32'h0;
      Register_inst43 <= 32'h0;
      Register_inst44 <= 32'h0;
      Register_inst45 <= 32'h0;
      Register_inst46 <= 32'h0;
      Register_inst47 <= 32'h0;
      Register_inst48 <= 32'h0;
      Register_inst49 <= 32'h0;
      Register_inst50 <= 32'h0;
      Register_inst51 <= 32'h0;
      Register_inst52 <= 32'h0;
      Register_inst53 <= 32'h0;
      Register_inst54 <= 32'h0;
      Register_inst55 <= 32'h0;
      Register_inst56 <= 32'h0;
      Register_inst57 <= 32'h0;
      Register_inst58 <= 32'h0;
      Register_inst59 <= 32'h0;
      Register_inst60 <= 32'h0;
      Register_inst61 <= 32'h0;
      Register_inst62 <= 32'h0;
      Register_inst63 <= 32'h0;
      Register_inst64 <= 32'h0;
      Register_inst65 <= 32'h0;
      Register_inst66 <= 32'h0;
      Register_inst67 <= 32'h0;
      Register_inst68 <= 32'h0;
      Register_inst69 <= 32'h0;
      Register_inst70 <= 32'h0;
      Register_inst71 <= 32'h0;
      Register_inst72 <= 32'h0;
      Register_inst73 <= 32'h0;
      Register_inst74 <= 32'h0;
      Register_inst75 <= 32'h0;
      Register_inst76 <= 32'h0;
      Register_inst77 <= 32'h0;
      Register_inst78 <= 32'h0;
      Register_inst79 <= 32'h0;
      Register_inst80 <= 32'h0;
      Register_inst81 <= 32'h0;
      Register_inst82 <= 32'h0;
      Register_inst83 <= 32'h0;
      Register_inst84 <= 32'h0;
      Register_inst85 <= 32'h0;
      Register_inst86 <= 32'h0;
      Register_inst87 <= 32'h0;
      Register_inst88 <= 32'h0;
      Register_inst89 <= 32'h0;
      Register_inst90 <= 32'h0;
      Register_inst91 <= 32'h0;
      Register_inst92 <= 32'h0;
      Register_inst93 <= 32'h0;
      Register_inst94 <= 32'h0;
      Register_inst95 <= 32'h0;
      Register_inst96 <= 32'h0;
      Register_inst97 <= 32'h0;
      Register_inst98 <= 32'h0;
      Register_inst99 <= 32'h0;
      Register_inst100 <= 32'h0;
      Register_inst101 <= 32'h0;
      Register_inst102 <= 32'h0;
      Register_inst103 <= 32'h0;
      Register_inst104 <= 32'h0;
      Register_inst105 <= 32'h0;
      Register_inst106 <= 32'h0;
      Register_inst107 <= 32'h0;
      Register_inst108 <= 32'h0;
      Register_inst109 <= 32'h0;
      Register_inst110 <= 32'h0;
      Register_inst111 <= 32'h0;
      Register_inst112 <= 32'h0;
      Register_inst113 <= 32'h0;
      Register_inst114 <= 32'h0;
      Register_inst115 <= 32'h0;
      Register_inst116 <= 32'h0;
      Register_inst117 <= 32'h0;
      Register_inst118 <= 32'h0;
      Register_inst119 <= 32'h0;
      Register_inst120 <= 32'h0;
      Register_inst121 <= 32'h0;
      Register_inst122 <= 32'h0;
      Register_inst123 <= 32'h0;
      Register_inst124 <= 32'h0;
      Register_inst125 <= 32'h0;
      Register_inst126 <= 32'h0;
      Register_inst127 <= 32'h0;
      Register_inst128 <= 32'h0;
      Register_inst129 <= 32'h0;
      Register_inst130 <= 32'h0;
      Register_inst131 <= 32'h0;
      Register_inst132 <= 32'h0;
      Register_inst133 <= 32'h0;
      Register_inst134 <= 32'h0;
      Register_inst135 <= 32'h0;
      Register_inst136 <= 32'h0;
      Register_inst137 <= 32'h0;
      Register_inst138 <= 32'h0;
      Register_inst139 <= 32'h0;
      Register_inst140 <= 32'h0;
      Register_inst141 <= 32'h0;
      Register_inst142 <= 32'h0;
      Register_inst143 <= 32'h0;
      Register_inst144 <= 32'h0;
      Register_inst145 <= 32'h0;
      Register_inst146 <= 32'h0;
      Register_inst147 <= 32'h0;
      Register_inst148 <= 32'h0;
      Register_inst149 <= 32'h0;
      Register_inst150 <= 32'h0;
      Register_inst151 <= 32'h0;
      Register_inst152 <= 32'h0;
      Register_inst153 <= 32'h0;
      Register_inst154 <= 32'h0;
      Register_inst155 <= 32'h0;
      Register_inst156 <= 32'h0;
      Register_inst157 <= 32'h0;
      Register_inst158 <= 32'h0;
      Register_inst159 <= 32'h0;
      Register_inst160 <= 32'h0;
      Register_inst161 <= 32'h0;
      Register_inst162 <= 32'h0;
      Register_inst163 <= 32'h0;
      Register_inst164 <= 32'h0;
      Register_inst165 <= 32'h0;
      Register_inst166 <= 32'h0;
      Register_inst167 <= 32'h0;
      Register_inst168 <= 32'h0;
      Register_inst169 <= 32'h0;
      Register_inst170 <= 32'h0;
      Register_inst171 <= 32'h0;
      Register_inst172 <= 32'h0;
      Register_inst173 <= 32'h0;
      Register_inst174 <= 32'h0;
      Register_inst175 <= 32'h0;
      Register_inst176 <= 32'h0;
      Register_inst177 <= 32'h0;
      Register_inst178 <= 32'h0;
      Register_inst179 <= 32'h0;
      Register_inst180 <= 32'h0;
      Register_inst181 <= 32'h0;
      Register_inst182 <= 32'h0;
      Register_inst183 <= 32'h0;
      Register_inst184 <= 32'h0;
      Register_inst185 <= 32'h0;
      Register_inst186 <= 32'h0;
      Register_inst187 <= 32'h0;
      Register_inst188 <= 32'h0;
      Register_inst189 <= 32'h0;
      Register_inst190 <= 32'h0;
      Register_inst191 <= 32'h0;
      Register_inst192 <= 32'h0;
      Register_inst193 <= 32'h0;
      Register_inst194 <= 32'h0;
      Register_inst195 <= 32'h0;
      Register_inst196 <= 32'h0;
      Register_inst197 <= 32'h0;
      Register_inst198 <= 32'h0;
      Register_inst199 <= 32'h0;
      Register_inst200 <= 32'h0;
      Register_inst201 <= 32'h0;
      Register_inst202 <= 32'h0;
      Register_inst203 <= 32'h0;
      Register_inst204 <= 32'h0;
      Register_inst205 <= 32'h0;
      Register_inst206 <= 32'h0;
      Register_inst207 <= 32'h0;
      Register_inst208 <= 32'h0;
      Register_inst209 <= 32'h0;
      Register_inst210 <= 32'h0;
      Register_inst211 <= 32'h0;
      Register_inst212 <= 32'h0;
      Register_inst213 <= 32'h0;
      Register_inst214 <= 32'h0;
      Register_inst215 <= 32'h0;
      Register_inst216 <= 32'h0;
      Register_inst217 <= 32'h0;
      Register_inst218 <= 32'h0;
      Register_inst219 <= 32'h0;
      Register_inst220 <= 32'h0;
      Register_inst221 <= 32'h0;
      Register_inst222 <= 32'h0;
      Register_inst223 <= 32'h0;
      Register_inst224 <= 32'h0;
      Register_inst225 <= 32'h0;
      Register_inst226 <= 32'h0;
      Register_inst227 <= 32'h0;
      Register_inst228 <= 32'h0;
      Register_inst229 <= 32'h0;
      Register_inst230 <= 32'h0;
      Register_inst231 <= 32'h0;
      Register_inst232 <= 32'h0;
      Register_inst233 <= 32'h0;
      Register_inst234 <= 32'h0;
      Register_inst235 <= 32'h0;
      Register_inst236 <= 32'h0;
      Register_inst237 <= 32'h0;
      Register_inst238 <= 32'h0;
      Register_inst239 <= 32'h0;
      Register_inst240 <= 32'h0;
      Register_inst241 <= 32'h0;
      Register_inst242 <= 32'h0;
      Register_inst243 <= 32'h0;
      Register_inst244 <= 32'h0;
      Register_inst245 <= 32'h0;
      Register_inst246 <= 32'h0;
      Register_inst247 <= 32'h0;
      Register_inst248 <= 32'h0;
      Register_inst249 <= 32'h0;
      Register_inst250 <= 32'h0;
      Register_inst251 <= 32'h0;
      Register_inst252 <= 32'h0;
      Register_inst253 <= 32'h0;
      Register_inst254 <= 32'h0;
      Register_inst255 <= 32'h0;
    end
    else begin
      automatic logic [31:0]      _T_0 = write_0.data;
      automatic logic [7:0]       _T_1 = write_0.addr;
      automatic logic [1:0][31:0] _T_2 = {{Register_inst0}, {_T_0}};
      automatic logic [1:0][31:0] _T_3 = {{Register_inst1}, {_T_0}};
      automatic logic [1:0][31:0] _T_4 = {{Register_inst2}, {_T_0}};
      automatic logic [1:0][31:0] _T_5 = {{Register_inst3}, {_T_0}};
      automatic logic [1:0][31:0] _T_6 = {{Register_inst4}, {_T_0}};
      automatic logic [1:0][31:0] _T_7 = {{Register_inst5}, {_T_0}};
      automatic logic [1:0][31:0] _T_8 = {{Register_inst6}, {_T_0}};
      automatic logic [1:0][31:0] _T_9 = {{Register_inst7}, {_T_0}};
      automatic logic [1:0][31:0] _T_10 = {{Register_inst8}, {_T_0}};
      automatic logic [1:0][31:0] _T_11 = {{Register_inst9}, {_T_0}};
      automatic logic [1:0][31:0] _T_12 = {{Register_inst10}, {_T_0}};
      automatic logic [1:0][31:0] _T_13 = {{Register_inst11}, {_T_0}};
      automatic logic [1:0][31:0] _T_14 = {{Register_inst12}, {_T_0}};
      automatic logic [1:0][31:0] _T_15 = {{Register_inst13}, {_T_0}};
      automatic logic [1:0][31:0] _T_16 = {{Register_inst14}, {_T_0}};
      automatic logic [1:0][31:0] _T_17 = {{Register_inst15}, {_T_0}};
      automatic logic [1:0][31:0] _T_18 = {{Register_inst16}, {_T_0}};
      automatic logic [1:0][31:0] _T_19 = {{Register_inst17}, {_T_0}};
      automatic logic [1:0][31:0] _T_20 = {{Register_inst18}, {_T_0}};
      automatic logic [1:0][31:0] _T_21 = {{Register_inst19}, {_T_0}};
      automatic logic [1:0][31:0] _T_22 = {{Register_inst20}, {_T_0}};
      automatic logic [1:0][31:0] _T_23 = {{Register_inst21}, {_T_0}};
      automatic logic [1:0][31:0] _T_24 = {{Register_inst22}, {_T_0}};
      automatic logic [1:0][31:0] _T_25 = {{Register_inst23}, {_T_0}};
      automatic logic [1:0][31:0] _T_26 = {{Register_inst24}, {_T_0}};
      automatic logic [1:0][31:0] _T_27 = {{Register_inst25}, {_T_0}};
      automatic logic [1:0][31:0] _T_28 = {{Register_inst26}, {_T_0}};
      automatic logic [1:0][31:0] _T_29 = {{Register_inst27}, {_T_0}};
      automatic logic [1:0][31:0] _T_30 = {{Register_inst28}, {_T_0}};
      automatic logic [1:0][31:0] _T_31 = {{Register_inst29}, {_T_0}};
      automatic logic [1:0][31:0] _T_32 = {{Register_inst30}, {_T_0}};
      automatic logic [1:0][31:0] _T_33 = {{Register_inst31}, {_T_0}};
      automatic logic [1:0][31:0] _T_34 = {{Register_inst32}, {_T_0}};
      automatic logic [1:0][31:0] _T_35 = {{Register_inst33}, {_T_0}};
      automatic logic [1:0][31:0] _T_36 = {{Register_inst34}, {_T_0}};
      automatic logic [1:0][31:0] _T_37 = {{Register_inst35}, {_T_0}};
      automatic logic [1:0][31:0] _T_38 = {{Register_inst36}, {_T_0}};
      automatic logic [1:0][31:0] _T_39 = {{Register_inst37}, {_T_0}};
      automatic logic [1:0][31:0] _T_40 = {{Register_inst38}, {_T_0}};
      automatic logic [1:0][31:0] _T_41 = {{Register_inst39}, {_T_0}};
      automatic logic [1:0][31:0] _T_42 = {{Register_inst40}, {_T_0}};
      automatic logic [1:0][31:0] _T_43 = {{Register_inst41}, {_T_0}};
      automatic logic [1:0][31:0] _T_44 = {{Register_inst42}, {_T_0}};
      automatic logic [1:0][31:0] _T_45 = {{Register_inst43}, {_T_0}};
      automatic logic [1:0][31:0] _T_46 = {{Register_inst44}, {_T_0}};
      automatic logic [1:0][31:0] _T_47 = {{Register_inst45}, {_T_0}};
      automatic logic [1:0][31:0] _T_48 = {{Register_inst46}, {_T_0}};
      automatic logic [1:0][31:0] _T_49 = {{Register_inst47}, {_T_0}};
      automatic logic [1:0][31:0] _T_50 = {{Register_inst48}, {_T_0}};
      automatic logic [1:0][31:0] _T_51 = {{Register_inst49}, {_T_0}};
      automatic logic [1:0][31:0] _T_52 = {{Register_inst50}, {_T_0}};
      automatic logic [1:0][31:0] _T_53 = {{Register_inst51}, {_T_0}};
      automatic logic [1:0][31:0] _T_54 = {{Register_inst52}, {_T_0}};
      automatic logic [1:0][31:0] _T_55 = {{Register_inst53}, {_T_0}};
      automatic logic [1:0][31:0] _T_56 = {{Register_inst54}, {_T_0}};
      automatic logic [1:0][31:0] _T_57 = {{Register_inst55}, {_T_0}};
      automatic logic [1:0][31:0] _T_58 = {{Register_inst56}, {_T_0}};
      automatic logic [1:0][31:0] _T_59 = {{Register_inst57}, {_T_0}};
      automatic logic [1:0][31:0] _T_60 = {{Register_inst58}, {_T_0}};
      automatic logic [1:0][31:0] _T_61 = {{Register_inst59}, {_T_0}};
      automatic logic [1:0][31:0] _T_62 = {{Register_inst60}, {_T_0}};
      automatic logic [1:0][31:0] _T_63 = {{Register_inst61}, {_T_0}};
      automatic logic [1:0][31:0] _T_64 = {{Register_inst62}, {_T_0}};
      automatic logic [1:0][31:0] _T_65 = {{Register_inst63}, {_T_0}};
      automatic logic [1:0][31:0] _T_66 = {{Register_inst64}, {_T_0}};
      automatic logic [1:0][31:0] _T_67 = {{Register_inst65}, {_T_0}};
      automatic logic [1:0][31:0] _T_68 = {{Register_inst66}, {_T_0}};
      automatic logic [1:0][31:0] _T_69 = {{Register_inst67}, {_T_0}};
      automatic logic [1:0][31:0] _T_70 = {{Register_inst68}, {_T_0}};
      automatic logic [1:0][31:0] _T_71 = {{Register_inst69}, {_T_0}};
      automatic logic [1:0][31:0] _T_72 = {{Register_inst70}, {_T_0}};
      automatic logic [1:0][31:0] _T_73 = {{Register_inst71}, {_T_0}};
      automatic logic [1:0][31:0] _T_74 = {{Register_inst72}, {_T_0}};
      automatic logic [1:0][31:0] _T_75 = {{Register_inst73}, {_T_0}};
      automatic logic [1:0][31:0] _T_76 = {{Register_inst74}, {_T_0}};
      automatic logic [1:0][31:0] _T_77 = {{Register_inst75}, {_T_0}};
      automatic logic [1:0][31:0] _T_78 = {{Register_inst76}, {_T_0}};
      automatic logic [1:0][31:0] _T_79 = {{Register_inst77}, {_T_0}};
      automatic logic [1:0][31:0] _T_80 = {{Register_inst78}, {_T_0}};
      automatic logic [1:0][31:0] _T_81 = {{Register_inst79}, {_T_0}};
      automatic logic [1:0][31:0] _T_82 = {{Register_inst80}, {_T_0}};
      automatic logic [1:0][31:0] _T_83 = {{Register_inst81}, {_T_0}};
      automatic logic [1:0][31:0] _T_84 = {{Register_inst82}, {_T_0}};
      automatic logic [1:0][31:0] _T_85 = {{Register_inst83}, {_T_0}};
      automatic logic [1:0][31:0] _T_86 = {{Register_inst84}, {_T_0}};
      automatic logic [1:0][31:0] _T_87 = {{Register_inst85}, {_T_0}};
      automatic logic [1:0][31:0] _T_88 = {{Register_inst86}, {_T_0}};
      automatic logic [1:0][31:0] _T_89 = {{Register_inst87}, {_T_0}};
      automatic logic [1:0][31:0] _T_90 = {{Register_inst88}, {_T_0}};
      automatic logic [1:0][31:0] _T_91 = {{Register_inst89}, {_T_0}};
      automatic logic [1:0][31:0] _T_92 = {{Register_inst90}, {_T_0}};
      automatic logic [1:0][31:0] _T_93 = {{Register_inst91}, {_T_0}};
      automatic logic [1:0][31:0] _T_94 = {{Register_inst92}, {_T_0}};
      automatic logic [1:0][31:0] _T_95 = {{Register_inst93}, {_T_0}};
      automatic logic [1:0][31:0] _T_96 = {{Register_inst94}, {_T_0}};
      automatic logic [1:0][31:0] _T_97 = {{Register_inst95}, {_T_0}};
      automatic logic [1:0][31:0] _T_98 = {{Register_inst96}, {_T_0}};
      automatic logic [1:0][31:0] _T_99 = {{Register_inst97}, {_T_0}};
      automatic logic [1:0][31:0] _T_100 = {{Register_inst98}, {_T_0}};
      automatic logic [1:0][31:0] _T_101 = {{Register_inst99}, {_T_0}};
      automatic logic [1:0][31:0] _T_102 = {{Register_inst100}, {_T_0}};
      automatic logic [1:0][31:0] _T_103 = {{Register_inst101}, {_T_0}};
      automatic logic [1:0][31:0] _T_104 = {{Register_inst102}, {_T_0}};
      automatic logic [1:0][31:0] _T_105 = {{Register_inst103}, {_T_0}};
      automatic logic [1:0][31:0] _T_106 = {{Register_inst104}, {_T_0}};
      automatic logic [1:0][31:0] _T_107 = {{Register_inst105}, {_T_0}};
      automatic logic [1:0][31:0] _T_108 = {{Register_inst106}, {_T_0}};
      automatic logic [1:0][31:0] _T_109 = {{Register_inst107}, {_T_0}};
      automatic logic [1:0][31:0] _T_110 = {{Register_inst108}, {_T_0}};
      automatic logic [1:0][31:0] _T_111 = {{Register_inst109}, {_T_0}};
      automatic logic [1:0][31:0] _T_112 = {{Register_inst110}, {_T_0}};
      automatic logic [1:0][31:0] _T_113 = {{Register_inst111}, {_T_0}};
      automatic logic [1:0][31:0] _T_114 = {{Register_inst112}, {_T_0}};
      automatic logic [1:0][31:0] _T_115 = {{Register_inst113}, {_T_0}};
      automatic logic [1:0][31:0] _T_116 = {{Register_inst114}, {_T_0}};
      automatic logic [1:0][31:0] _T_117 = {{Register_inst115}, {_T_0}};
      automatic logic [1:0][31:0] _T_118 = {{Register_inst116}, {_T_0}};
      automatic logic [1:0][31:0] _T_119 = {{Register_inst117}, {_T_0}};
      automatic logic [1:0][31:0] _T_120 = {{Register_inst118}, {_T_0}};
      automatic logic [1:0][31:0] _T_121 = {{Register_inst119}, {_T_0}};
      automatic logic [1:0][31:0] _T_122 = {{Register_inst120}, {_T_0}};
      automatic logic [1:0][31:0] _T_123 = {{Register_inst121}, {_T_0}};
      automatic logic [1:0][31:0] _T_124 = {{Register_inst122}, {_T_0}};
      automatic logic [1:0][31:0] _T_125 = {{Register_inst123}, {_T_0}};
      automatic logic [1:0][31:0] _T_126 = {{Register_inst124}, {_T_0}};
      automatic logic [1:0][31:0] _T_127 = {{Register_inst125}, {_T_0}};
      automatic logic [1:0][31:0] _T_128 = {{Register_inst126}, {_T_0}};
      automatic logic [1:0][31:0] _T_129 = {{Register_inst127}, {_T_0}};
      automatic logic [1:0][31:0] _T_130 = {{Register_inst128}, {_T_0}};
      automatic logic [1:0][31:0] _T_131 = {{Register_inst129}, {_T_0}};
      automatic logic [1:0][31:0] _T_132 = {{Register_inst130}, {_T_0}};
      automatic logic [1:0][31:0] _T_133 = {{Register_inst131}, {_T_0}};
      automatic logic [1:0][31:0] _T_134 = {{Register_inst132}, {_T_0}};
      automatic logic [1:0][31:0] _T_135 = {{Register_inst133}, {_T_0}};
      automatic logic [1:0][31:0] _T_136 = {{Register_inst134}, {_T_0}};
      automatic logic [1:0][31:0] _T_137 = {{Register_inst135}, {_T_0}};
      automatic logic [1:0][31:0] _T_138 = {{Register_inst136}, {_T_0}};
      automatic logic [1:0][31:0] _T_139 = {{Register_inst137}, {_T_0}};
      automatic logic [1:0][31:0] _T_140 = {{Register_inst138}, {_T_0}};
      automatic logic [1:0][31:0] _T_141 = {{Register_inst139}, {_T_0}};
      automatic logic [1:0][31:0] _T_142 = {{Register_inst140}, {_T_0}};
      automatic logic [1:0][31:0] _T_143 = {{Register_inst141}, {_T_0}};
      automatic logic [1:0][31:0] _T_144 = {{Register_inst142}, {_T_0}};
      automatic logic [1:0][31:0] _T_145 = {{Register_inst143}, {_T_0}};
      automatic logic [1:0][31:0] _T_146 = {{Register_inst144}, {_T_0}};
      automatic logic [1:0][31:0] _T_147 = {{Register_inst145}, {_T_0}};
      automatic logic [1:0][31:0] _T_148 = {{Register_inst146}, {_T_0}};
      automatic logic [1:0][31:0] _T_149 = {{Register_inst147}, {_T_0}};
      automatic logic [1:0][31:0] _T_150 = {{Register_inst148}, {_T_0}};
      automatic logic [1:0][31:0] _T_151 = {{Register_inst149}, {_T_0}};
      automatic logic [1:0][31:0] _T_152 = {{Register_inst150}, {_T_0}};
      automatic logic [1:0][31:0] _T_153 = {{Register_inst151}, {_T_0}};
      automatic logic [1:0][31:0] _T_154 = {{Register_inst152}, {_T_0}};
      automatic logic [1:0][31:0] _T_155 = {{Register_inst153}, {_T_0}};
      automatic logic [1:0][31:0] _T_156 = {{Register_inst154}, {_T_0}};
      automatic logic [1:0][31:0] _T_157 = {{Register_inst155}, {_T_0}};
      automatic logic [1:0][31:0] _T_158 = {{Register_inst156}, {_T_0}};
      automatic logic [1:0][31:0] _T_159 = {{Register_inst157}, {_T_0}};
      automatic logic [1:0][31:0] _T_160 = {{Register_inst158}, {_T_0}};
      automatic logic [1:0][31:0] _T_161 = {{Register_inst159}, {_T_0}};
      automatic logic [1:0][31:0] _T_162 = {{Register_inst160}, {_T_0}};
      automatic logic [1:0][31:0] _T_163 = {{Register_inst161}, {_T_0}};
      automatic logic [1:0][31:0] _T_164 = {{Register_inst162}, {_T_0}};
      automatic logic [1:0][31:0] _T_165 = {{Register_inst163}, {_T_0}};
      automatic logic [1:0][31:0] _T_166 = {{Register_inst164}, {_T_0}};
      automatic logic [1:0][31:0] _T_167 = {{Register_inst165}, {_T_0}};
      automatic logic [1:0][31:0] _T_168 = {{Register_inst166}, {_T_0}};
      automatic logic [1:0][31:0] _T_169 = {{Register_inst167}, {_T_0}};
      automatic logic [1:0][31:0] _T_170 = {{Register_inst168}, {_T_0}};
      automatic logic [1:0][31:0] _T_171 = {{Register_inst169}, {_T_0}};
      automatic logic [1:0][31:0] _T_172 = {{Register_inst170}, {_T_0}};
      automatic logic [1:0][31:0] _T_173 = {{Register_inst171}, {_T_0}};
      automatic logic [1:0][31:0] _T_174 = {{Register_inst172}, {_T_0}};
      automatic logic [1:0][31:0] _T_175 = {{Register_inst173}, {_T_0}};
      automatic logic [1:0][31:0] _T_176 = {{Register_inst174}, {_T_0}};
      automatic logic [1:0][31:0] _T_177 = {{Register_inst175}, {_T_0}};
      automatic logic [1:0][31:0] _T_178 = {{Register_inst176}, {_T_0}};
      automatic logic [1:0][31:0] _T_179 = {{Register_inst177}, {_T_0}};
      automatic logic [1:0][31:0] _T_180 = {{Register_inst178}, {_T_0}};
      automatic logic [1:0][31:0] _T_181 = {{Register_inst179}, {_T_0}};
      automatic logic [1:0][31:0] _T_182 = {{Register_inst180}, {_T_0}};
      automatic logic [1:0][31:0] _T_183 = {{Register_inst181}, {_T_0}};
      automatic logic [1:0][31:0] _T_184 = {{Register_inst182}, {_T_0}};
      automatic logic [1:0][31:0] _T_185 = {{Register_inst183}, {_T_0}};
      automatic logic [1:0][31:0] _T_186 = {{Register_inst184}, {_T_0}};
      automatic logic [1:0][31:0] _T_187 = {{Register_inst185}, {_T_0}};
      automatic logic [1:0][31:0] _T_188 = {{Register_inst186}, {_T_0}};
      automatic logic [1:0][31:0] _T_189 = {{Register_inst187}, {_T_0}};
      automatic logic [1:0][31:0] _T_190 = {{Register_inst188}, {_T_0}};
      automatic logic [1:0][31:0] _T_191 = {{Register_inst189}, {_T_0}};
      automatic logic [1:0][31:0] _T_192 = {{Register_inst190}, {_T_0}};
      automatic logic [1:0][31:0] _T_193 = {{Register_inst191}, {_T_0}};
      automatic logic [1:0][31:0] _T_194 = {{Register_inst192}, {_T_0}};
      automatic logic [1:0][31:0] _T_195 = {{Register_inst193}, {_T_0}};
      automatic logic [1:0][31:0] _T_196 = {{Register_inst194}, {_T_0}};
      automatic logic [1:0][31:0] _T_197 = {{Register_inst195}, {_T_0}};
      automatic logic [1:0][31:0] _T_198 = {{Register_inst196}, {_T_0}};
      automatic logic [1:0][31:0] _T_199 = {{Register_inst197}, {_T_0}};
      automatic logic [1:0][31:0] _T_200 = {{Register_inst198}, {_T_0}};
      automatic logic [1:0][31:0] _T_201 = {{Register_inst199}, {_T_0}};
      automatic logic [1:0][31:0] _T_202 = {{Register_inst200}, {_T_0}};
      automatic logic [1:0][31:0] _T_203 = {{Register_inst201}, {_T_0}};
      automatic logic [1:0][31:0] _T_204 = {{Register_inst202}, {_T_0}};
      automatic logic [1:0][31:0] _T_205 = {{Register_inst203}, {_T_0}};
      automatic logic [1:0][31:0] _T_206 = {{Register_inst204}, {_T_0}};
      automatic logic [1:0][31:0] _T_207 = {{Register_inst205}, {_T_0}};
      automatic logic [1:0][31:0] _T_208 = {{Register_inst206}, {_T_0}};
      automatic logic [1:0][31:0] _T_209 = {{Register_inst207}, {_T_0}};
      automatic logic [1:0][31:0] _T_210 = {{Register_inst208}, {_T_0}};
      automatic logic [1:0][31:0] _T_211 = {{Register_inst209}, {_T_0}};
      automatic logic [1:0][31:0] _T_212 = {{Register_inst210}, {_T_0}};
      automatic logic [1:0][31:0] _T_213 = {{Register_inst211}, {_T_0}};
      automatic logic [1:0][31:0] _T_214 = {{Register_inst212}, {_T_0}};
      automatic logic [1:0][31:0] _T_215 = {{Register_inst213}, {_T_0}};
      automatic logic [1:0][31:0] _T_216 = {{Register_inst214}, {_T_0}};
      automatic logic [1:0][31:0] _T_217 = {{Register_inst215}, {_T_0}};
      automatic logic [1:0][31:0] _T_218 = {{Register_inst216}, {_T_0}};
      automatic logic [1:0][31:0] _T_219 = {{Register_inst217}, {_T_0}};
      automatic logic [1:0][31:0] _T_220 = {{Register_inst218}, {_T_0}};
      automatic logic [1:0][31:0] _T_221 = {{Register_inst219}, {_T_0}};
      automatic logic [1:0][31:0] _T_222 = {{Register_inst220}, {_T_0}};
      automatic logic [1:0][31:0] _T_223 = {{Register_inst221}, {_T_0}};
      automatic logic [1:0][31:0] _T_224 = {{Register_inst222}, {_T_0}};
      automatic logic [1:0][31:0] _T_225 = {{Register_inst223}, {_T_0}};
      automatic logic [1:0][31:0] _T_226 = {{Register_inst224}, {_T_0}};
      automatic logic [1:0][31:0] _T_227 = {{Register_inst225}, {_T_0}};
      automatic logic [1:0][31:0] _T_228 = {{Register_inst226}, {_T_0}};
      automatic logic [1:0][31:0] _T_229 = {{Register_inst227}, {_T_0}};
      automatic logic [1:0][31:0] _T_230 = {{Register_inst228}, {_T_0}};
      automatic logic [1:0][31:0] _T_231 = {{Register_inst229}, {_T_0}};
      automatic logic [1:0][31:0] _T_232 = {{Register_inst230}, {_T_0}};
      automatic logic [1:0][31:0] _T_233 = {{Register_inst231}, {_T_0}};
      automatic logic [1:0][31:0] _T_234 = {{Register_inst232}, {_T_0}};
      automatic logic [1:0][31:0] _T_235 = {{Register_inst233}, {_T_0}};
      automatic logic [1:0][31:0] _T_236 = {{Register_inst234}, {_T_0}};
      automatic logic [1:0][31:0] _T_237 = {{Register_inst235}, {_T_0}};
      automatic logic [1:0][31:0] _T_238 = {{Register_inst236}, {_T_0}};
      automatic logic [1:0][31:0] _T_239 = {{Register_inst237}, {_T_0}};
      automatic logic [1:0][31:0] _T_240 = {{Register_inst238}, {_T_0}};
      automatic logic [1:0][31:0] _T_241 = {{Register_inst239}, {_T_0}};
      automatic logic [1:0][31:0] _T_242 = {{Register_inst240}, {_T_0}};
      automatic logic [1:0][31:0] _T_243 = {{Register_inst241}, {_T_0}};
      automatic logic [1:0][31:0] _T_244 = {{Register_inst242}, {_T_0}};
      automatic logic [1:0][31:0] _T_245 = {{Register_inst243}, {_T_0}};
      automatic logic [1:0][31:0] _T_246 = {{Register_inst244}, {_T_0}};
      automatic logic [1:0][31:0] _T_247 = {{Register_inst245}, {_T_0}};
      automatic logic [1:0][31:0] _T_248 = {{Register_inst246}, {_T_0}};
      automatic logic [1:0][31:0] _T_249 = {{Register_inst247}, {_T_0}};
      automatic logic [1:0][31:0] _T_250 = {{Register_inst248}, {_T_0}};
      automatic logic [1:0][31:0] _T_251 = {{Register_inst249}, {_T_0}};
      automatic logic [1:0][31:0] _T_252 = {{Register_inst250}, {_T_0}};
      automatic logic [1:0][31:0] _T_253 = {{Register_inst251}, {_T_0}};
      automatic logic [1:0][31:0] _T_254 = {{Register_inst252}, {_T_0}};
      automatic logic [1:0][31:0] _T_255 = {{Register_inst253}, {_T_0}};
      automatic logic [1:0][31:0] _T_256 = {{Register_inst254}, {_T_0}};
      automatic logic [1:0][31:0] _T_257 = {{Register_inst255}, {_T_0}};

      Register_inst0 <= _T_2[_T_1 == 8'h0 & write_0_en];
      Register_inst1 <= _T_3[_T_1 == 8'h1 & write_0_en];
      Register_inst2 <= _T_4[_T_1 == 8'h2 & write_0_en];
      Register_inst3 <= _T_5[_T_1 == 8'h3 & write_0_en];
      Register_inst4 <= _T_6[_T_1 == 8'h4 & write_0_en];
      Register_inst5 <= _T_7[_T_1 == 8'h5 & write_0_en];
      Register_inst6 <= _T_8[_T_1 == 8'h6 & write_0_en];
      Register_inst7 <= _T_9[_T_1 == 8'h7 & write_0_en];
      Register_inst8 <= _T_10[_T_1 == 8'h8 & write_0_en];
      Register_inst9 <= _T_11[_T_1 == 8'h9 & write_0_en];
      Register_inst10 <= _T_12[_T_1 == 8'hA & write_0_en];
      Register_inst11 <= _T_13[_T_1 == 8'hB & write_0_en];
      Register_inst12 <= _T_14[_T_1 == 8'hC & write_0_en];
      Register_inst13 <= _T_15[_T_1 == 8'hD & write_0_en];
      Register_inst14 <= _T_16[_T_1 == 8'hE & write_0_en];
      Register_inst15 <= _T_17[_T_1 == 8'hF & write_0_en];
      Register_inst16 <= _T_18[_T_1 == 8'h10 & write_0_en];
      Register_inst17 <= _T_19[_T_1 == 8'h11 & write_0_en];
      Register_inst18 <= _T_20[_T_1 == 8'h12 & write_0_en];
      Register_inst19 <= _T_21[_T_1 == 8'h13 & write_0_en];
      Register_inst20 <= _T_22[_T_1 == 8'h14 & write_0_en];
      Register_inst21 <= _T_23[_T_1 == 8'h15 & write_0_en];
      Register_inst22 <= _T_24[_T_1 == 8'h16 & write_0_en];
      Register_inst23 <= _T_25[_T_1 == 8'h17 & write_0_en];
      Register_inst24 <= _T_26[_T_1 == 8'h18 & write_0_en];
      Register_inst25 <= _T_27[_T_1 == 8'h19 & write_0_en];
      Register_inst26 <= _T_28[_T_1 == 8'h1A & write_0_en];
      Register_inst27 <= _T_29[_T_1 == 8'h1B & write_0_en];
      Register_inst28 <= _T_30[_T_1 == 8'h1C & write_0_en];
      Register_inst29 <= _T_31[_T_1 == 8'h1D & write_0_en];
      Register_inst30 <= _T_32[_T_1 == 8'h1E & write_0_en];
      Register_inst31 <= _T_33[_T_1 == 8'h1F & write_0_en];
      Register_inst32 <= _T_34[_T_1 == 8'h20 & write_0_en];
      Register_inst33 <= _T_35[_T_1 == 8'h21 & write_0_en];
      Register_inst34 <= _T_36[_T_1 == 8'h22 & write_0_en];
      Register_inst35 <= _T_37[_T_1 == 8'h23 & write_0_en];
      Register_inst36 <= _T_38[_T_1 == 8'h24 & write_0_en];
      Register_inst37 <= _T_39[_T_1 == 8'h25 & write_0_en];
      Register_inst38 <= _T_40[_T_1 == 8'h26 & write_0_en];
      Register_inst39 <= _T_41[_T_1 == 8'h27 & write_0_en];
      Register_inst40 <= _T_42[_T_1 == 8'h28 & write_0_en];
      Register_inst41 <= _T_43[_T_1 == 8'h29 & write_0_en];
      Register_inst42 <= _T_44[_T_1 == 8'h2A & write_0_en];
      Register_inst43 <= _T_45[_T_1 == 8'h2B & write_0_en];
      Register_inst44 <= _T_46[_T_1 == 8'h2C & write_0_en];
      Register_inst45 <= _T_47[_T_1 == 8'h2D & write_0_en];
      Register_inst46 <= _T_48[_T_1 == 8'h2E & write_0_en];
      Register_inst47 <= _T_49[_T_1 == 8'h2F & write_0_en];
      Register_inst48 <= _T_50[_T_1 == 8'h30 & write_0_en];
      Register_inst49 <= _T_51[_T_1 == 8'h31 & write_0_en];
      Register_inst50 <= _T_52[_T_1 == 8'h32 & write_0_en];
      Register_inst51 <= _T_53[_T_1 == 8'h33 & write_0_en];
      Register_inst52 <= _T_54[_T_1 == 8'h34 & write_0_en];
      Register_inst53 <= _T_55[_T_1 == 8'h35 & write_0_en];
      Register_inst54 <= _T_56[_T_1 == 8'h36 & write_0_en];
      Register_inst55 <= _T_57[_T_1 == 8'h37 & write_0_en];
      Register_inst56 <= _T_58[_T_1 == 8'h38 & write_0_en];
      Register_inst57 <= _T_59[_T_1 == 8'h39 & write_0_en];
      Register_inst58 <= _T_60[_T_1 == 8'h3A & write_0_en];
      Register_inst59 <= _T_61[_T_1 == 8'h3B & write_0_en];
      Register_inst60 <= _T_62[_T_1 == 8'h3C & write_0_en];
      Register_inst61 <= _T_63[_T_1 == 8'h3D & write_0_en];
      Register_inst62 <= _T_64[_T_1 == 8'h3E & write_0_en];
      Register_inst63 <= _T_65[_T_1 == 8'h3F & write_0_en];
      Register_inst64 <= _T_66[_T_1 == 8'h40 & write_0_en];
      Register_inst65 <= _T_67[_T_1 == 8'h41 & write_0_en];
      Register_inst66 <= _T_68[_T_1 == 8'h42 & write_0_en];
      Register_inst67 <= _T_69[_T_1 == 8'h43 & write_0_en];
      Register_inst68 <= _T_70[_T_1 == 8'h44 & write_0_en];
      Register_inst69 <= _T_71[_T_1 == 8'h45 & write_0_en];
      Register_inst70 <= _T_72[_T_1 == 8'h46 & write_0_en];
      Register_inst71 <= _T_73[_T_1 == 8'h47 & write_0_en];
      Register_inst72 <= _T_74[_T_1 == 8'h48 & write_0_en];
      Register_inst73 <= _T_75[_T_1 == 8'h49 & write_0_en];
      Register_inst74 <= _T_76[_T_1 == 8'h4A & write_0_en];
      Register_inst75 <= _T_77[_T_1 == 8'h4B & write_0_en];
      Register_inst76 <= _T_78[_T_1 == 8'h4C & write_0_en];
      Register_inst77 <= _T_79[_T_1 == 8'h4D & write_0_en];
      Register_inst78 <= _T_80[_T_1 == 8'h4E & write_0_en];
      Register_inst79 <= _T_81[_T_1 == 8'h4F & write_0_en];
      Register_inst80 <= _T_82[_T_1 == 8'h50 & write_0_en];
      Register_inst81 <= _T_83[_T_1 == 8'h51 & write_0_en];
      Register_inst82 <= _T_84[_T_1 == 8'h52 & write_0_en];
      Register_inst83 <= _T_85[_T_1 == 8'h53 & write_0_en];
      Register_inst84 <= _T_86[_T_1 == 8'h54 & write_0_en];
      Register_inst85 <= _T_87[_T_1 == 8'h55 & write_0_en];
      Register_inst86 <= _T_88[_T_1 == 8'h56 & write_0_en];
      Register_inst87 <= _T_89[_T_1 == 8'h57 & write_0_en];
      Register_inst88 <= _T_90[_T_1 == 8'h58 & write_0_en];
      Register_inst89 <= _T_91[_T_1 == 8'h59 & write_0_en];
      Register_inst90 <= _T_92[_T_1 == 8'h5A & write_0_en];
      Register_inst91 <= _T_93[_T_1 == 8'h5B & write_0_en];
      Register_inst92 <= _T_94[_T_1 == 8'h5C & write_0_en];
      Register_inst93 <= _T_95[_T_1 == 8'h5D & write_0_en];
      Register_inst94 <= _T_96[_T_1 == 8'h5E & write_0_en];
      Register_inst95 <= _T_97[_T_1 == 8'h5F & write_0_en];
      Register_inst96 <= _T_98[_T_1 == 8'h60 & write_0_en];
      Register_inst97 <= _T_99[_T_1 == 8'h61 & write_0_en];
      Register_inst98 <= _T_100[_T_1 == 8'h62 & write_0_en];
      Register_inst99 <= _T_101[_T_1 == 8'h63 & write_0_en];
      Register_inst100 <= _T_102[_T_1 == 8'h64 & write_0_en];
      Register_inst101 <= _T_103[_T_1 == 8'h65 & write_0_en];
      Register_inst102 <= _T_104[_T_1 == 8'h66 & write_0_en];
      Register_inst103 <= _T_105[_T_1 == 8'h67 & write_0_en];
      Register_inst104 <= _T_106[_T_1 == 8'h68 & write_0_en];
      Register_inst105 <= _T_107[_T_1 == 8'h69 & write_0_en];
      Register_inst106 <= _T_108[_T_1 == 8'h6A & write_0_en];
      Register_inst107 <= _T_109[_T_1 == 8'h6B & write_0_en];
      Register_inst108 <= _T_110[_T_1 == 8'h6C & write_0_en];
      Register_inst109 <= _T_111[_T_1 == 8'h6D & write_0_en];
      Register_inst110 <= _T_112[_T_1 == 8'h6E & write_0_en];
      Register_inst111 <= _T_113[_T_1 == 8'h6F & write_0_en];
      Register_inst112 <= _T_114[_T_1 == 8'h70 & write_0_en];
      Register_inst113 <= _T_115[_T_1 == 8'h71 & write_0_en];
      Register_inst114 <= _T_116[_T_1 == 8'h72 & write_0_en];
      Register_inst115 <= _T_117[_T_1 == 8'h73 & write_0_en];
      Register_inst116 <= _T_118[_T_1 == 8'h74 & write_0_en];
      Register_inst117 <= _T_119[_T_1 == 8'h75 & write_0_en];
      Register_inst118 <= _T_120[_T_1 == 8'h76 & write_0_en];
      Register_inst119 <= _T_121[_T_1 == 8'h77 & write_0_en];
      Register_inst120 <= _T_122[_T_1 == 8'h78 & write_0_en];
      Register_inst121 <= _T_123[_T_1 == 8'h79 & write_0_en];
      Register_inst122 <= _T_124[_T_1 == 8'h7A & write_0_en];
      Register_inst123 <= _T_125[_T_1 == 8'h7B & write_0_en];
      Register_inst124 <= _T_126[_T_1 == 8'h7C & write_0_en];
      Register_inst125 <= _T_127[_T_1 == 8'h7D & write_0_en];
      Register_inst126 <= _T_128[_T_1 == 8'h7E & write_0_en];
      Register_inst127 <= _T_129[_T_1 == 8'h7F & write_0_en];
      Register_inst128 <= _T_130[_T_1 == 8'h80 & write_0_en];
      Register_inst129 <= _T_131[_T_1 == 8'h81 & write_0_en];
      Register_inst130 <= _T_132[_T_1 == 8'h82 & write_0_en];
      Register_inst131 <= _T_133[_T_1 == 8'h83 & write_0_en];
      Register_inst132 <= _T_134[_T_1 == 8'h84 & write_0_en];
      Register_inst133 <= _T_135[_T_1 == 8'h85 & write_0_en];
      Register_inst134 <= _T_136[_T_1 == 8'h86 & write_0_en];
      Register_inst135 <= _T_137[_T_1 == 8'h87 & write_0_en];
      Register_inst136 <= _T_138[_T_1 == 8'h88 & write_0_en];
      Register_inst137 <= _T_139[_T_1 == 8'h89 & write_0_en];
      Register_inst138 <= _T_140[_T_1 == 8'h8A & write_0_en];
      Register_inst139 <= _T_141[_T_1 == 8'h8B & write_0_en];
      Register_inst140 <= _T_142[_T_1 == 8'h8C & write_0_en];
      Register_inst141 <= _T_143[_T_1 == 8'h8D & write_0_en];
      Register_inst142 <= _T_144[_T_1 == 8'h8E & write_0_en];
      Register_inst143 <= _T_145[_T_1 == 8'h8F & write_0_en];
      Register_inst144 <= _T_146[_T_1 == 8'h90 & write_0_en];
      Register_inst145 <= _T_147[_T_1 == 8'h91 & write_0_en];
      Register_inst146 <= _T_148[_T_1 == 8'h92 & write_0_en];
      Register_inst147 <= _T_149[_T_1 == 8'h93 & write_0_en];
      Register_inst148 <= _T_150[_T_1 == 8'h94 & write_0_en];
      Register_inst149 <= _T_151[_T_1 == 8'h95 & write_0_en];
      Register_inst150 <= _T_152[_T_1 == 8'h96 & write_0_en];
      Register_inst151 <= _T_153[_T_1 == 8'h97 & write_0_en];
      Register_inst152 <= _T_154[_T_1 == 8'h98 & write_0_en];
      Register_inst153 <= _T_155[_T_1 == 8'h99 & write_0_en];
      Register_inst154 <= _T_156[_T_1 == 8'h9A & write_0_en];
      Register_inst155 <= _T_157[_T_1 == 8'h9B & write_0_en];
      Register_inst156 <= _T_158[_T_1 == 8'h9C & write_0_en];
      Register_inst157 <= _T_159[_T_1 == 8'h9D & write_0_en];
      Register_inst158 <= _T_160[_T_1 == 8'h9E & write_0_en];
      Register_inst159 <= _T_161[_T_1 == 8'h9F & write_0_en];
      Register_inst160 <= _T_162[_T_1 == 8'hA0 & write_0_en];
      Register_inst161 <= _T_163[_T_1 == 8'hA1 & write_0_en];
      Register_inst162 <= _T_164[_T_1 == 8'hA2 & write_0_en];
      Register_inst163 <= _T_165[_T_1 == 8'hA3 & write_0_en];
      Register_inst164 <= _T_166[_T_1 == 8'hA4 & write_0_en];
      Register_inst165 <= _T_167[_T_1 == 8'hA5 & write_0_en];
      Register_inst166 <= _T_168[_T_1 == 8'hA6 & write_0_en];
      Register_inst167 <= _T_169[_T_1 == 8'hA7 & write_0_en];
      Register_inst168 <= _T_170[_T_1 == 8'hA8 & write_0_en];
      Register_inst169 <= _T_171[_T_1 == 8'hA9 & write_0_en];
      Register_inst170 <= _T_172[_T_1 == 8'hAA & write_0_en];
      Register_inst171 <= _T_173[_T_1 == 8'hAB & write_0_en];
      Register_inst172 <= _T_174[_T_1 == 8'hAC & write_0_en];
      Register_inst173 <= _T_175[_T_1 == 8'hAD & write_0_en];
      Register_inst174 <= _T_176[_T_1 == 8'hAE & write_0_en];
      Register_inst175 <= _T_177[_T_1 == 8'hAF & write_0_en];
      Register_inst176 <= _T_178[_T_1 == 8'hB0 & write_0_en];
      Register_inst177 <= _T_179[_T_1 == 8'hB1 & write_0_en];
      Register_inst178 <= _T_180[_T_1 == 8'hB2 & write_0_en];
      Register_inst179 <= _T_181[_T_1 == 8'hB3 & write_0_en];
      Register_inst180 <= _T_182[_T_1 == 8'hB4 & write_0_en];
      Register_inst181 <= _T_183[_T_1 == 8'hB5 & write_0_en];
      Register_inst182 <= _T_184[_T_1 == 8'hB6 & write_0_en];
      Register_inst183 <= _T_185[_T_1 == 8'hB7 & write_0_en];
      Register_inst184 <= _T_186[_T_1 == 8'hB8 & write_0_en];
      Register_inst185 <= _T_187[_T_1 == 8'hB9 & write_0_en];
      Register_inst186 <= _T_188[_T_1 == 8'hBA & write_0_en];
      Register_inst187 <= _T_189[_T_1 == 8'hBB & write_0_en];
      Register_inst188 <= _T_190[_T_1 == 8'hBC & write_0_en];
      Register_inst189 <= _T_191[_T_1 == 8'hBD & write_0_en];
      Register_inst190 <= _T_192[_T_1 == 8'hBE & write_0_en];
      Register_inst191 <= _T_193[_T_1 == 8'hBF & write_0_en];
      Register_inst192 <= _T_194[_T_1 == 8'hC0 & write_0_en];
      Register_inst193 <= _T_195[_T_1 == 8'hC1 & write_0_en];
      Register_inst194 <= _T_196[_T_1 == 8'hC2 & write_0_en];
      Register_inst195 <= _T_197[_T_1 == 8'hC3 & write_0_en];
      Register_inst196 <= _T_198[_T_1 == 8'hC4 & write_0_en];
      Register_inst197 <= _T_199[_T_1 == 8'hC5 & write_0_en];
      Register_inst198 <= _T_200[_T_1 == 8'hC6 & write_0_en];
      Register_inst199 <= _T_201[_T_1 == 8'hC7 & write_0_en];
      Register_inst200 <= _T_202[_T_1 == 8'hC8 & write_0_en];
      Register_inst201 <= _T_203[_T_1 == 8'hC9 & write_0_en];
      Register_inst202 <= _T_204[_T_1 == 8'hCA & write_0_en];
      Register_inst203 <= _T_205[_T_1 == 8'hCB & write_0_en];
      Register_inst204 <= _T_206[_T_1 == 8'hCC & write_0_en];
      Register_inst205 <= _T_207[_T_1 == 8'hCD & write_0_en];
      Register_inst206 <= _T_208[_T_1 == 8'hCE & write_0_en];
      Register_inst207 <= _T_209[_T_1 == 8'hCF & write_0_en];
      Register_inst208 <= _T_210[_T_1 == 8'hD0 & write_0_en];
      Register_inst209 <= _T_211[_T_1 == 8'hD1 & write_0_en];
      Register_inst210 <= _T_212[_T_1 == 8'hD2 & write_0_en];
      Register_inst211 <= _T_213[_T_1 == 8'hD3 & write_0_en];
      Register_inst212 <= _T_214[_T_1 == 8'hD4 & write_0_en];
      Register_inst213 <= _T_215[_T_1 == 8'hD5 & write_0_en];
      Register_inst214 <= _T_216[_T_1 == 8'hD6 & write_0_en];
      Register_inst215 <= _T_217[_T_1 == 8'hD7 & write_0_en];
      Register_inst216 <= _T_218[_T_1 == 8'hD8 & write_0_en];
      Register_inst217 <= _T_219[_T_1 == 8'hD9 & write_0_en];
      Register_inst218 <= _T_220[_T_1 == 8'hDA & write_0_en];
      Register_inst219 <= _T_221[_T_1 == 8'hDB & write_0_en];
      Register_inst220 <= _T_222[_T_1 == 8'hDC & write_0_en];
      Register_inst221 <= _T_223[_T_1 == 8'hDD & write_0_en];
      Register_inst222 <= _T_224[_T_1 == 8'hDE & write_0_en];
      Register_inst223 <= _T_225[_T_1 == 8'hDF & write_0_en];
      Register_inst224 <= _T_226[_T_1 == 8'hE0 & write_0_en];
      Register_inst225 <= _T_227[_T_1 == 8'hE1 & write_0_en];
      Register_inst226 <= _T_228[_T_1 == 8'hE2 & write_0_en];
      Register_inst227 <= _T_229[_T_1 == 8'hE3 & write_0_en];
      Register_inst228 <= _T_230[_T_1 == 8'hE4 & write_0_en];
      Register_inst229 <= _T_231[_T_1 == 8'hE5 & write_0_en];
      Register_inst230 <= _T_232[_T_1 == 8'hE6 & write_0_en];
      Register_inst231 <= _T_233[_T_1 == 8'hE7 & write_0_en];
      Register_inst232 <= _T_234[_T_1 == 8'hE8 & write_0_en];
      Register_inst233 <= _T_235[_T_1 == 8'hE9 & write_0_en];
      Register_inst234 <= _T_236[_T_1 == 8'hEA & write_0_en];
      Register_inst235 <= _T_237[_T_1 == 8'hEB & write_0_en];
      Register_inst236 <= _T_238[_T_1 == 8'hEC & write_0_en];
      Register_inst237 <= _T_239[_T_1 == 8'hED & write_0_en];
      Register_inst238 <= _T_240[_T_1 == 8'hEE & write_0_en];
      Register_inst239 <= _T_241[_T_1 == 8'hEF & write_0_en];
      Register_inst240 <= _T_242[_T_1 == 8'hF0 & write_0_en];
      Register_inst241 <= _T_243[_T_1 == 8'hF1 & write_0_en];
      Register_inst242 <= _T_244[_T_1 == 8'hF2 & write_0_en];
      Register_inst243 <= _T_245[_T_1 == 8'hF3 & write_0_en];
      Register_inst244 <= _T_246[_T_1 == 8'hF4 & write_0_en];
      Register_inst245 <= _T_247[_T_1 == 8'hF5 & write_0_en];
      Register_inst246 <= _T_248[_T_1 == 8'hF6 & write_0_en];
      Register_inst247 <= _T_249[_T_1 == 8'hF7 & write_0_en];
      Register_inst248 <= _T_250[_T_1 == 8'hF8 & write_0_en];
      Register_inst249 <= _T_251[_T_1 == 8'hF9 & write_0_en];
      Register_inst250 <= _T_252[_T_1 == 8'hFA & write_0_en];
      Register_inst251 <= _T_253[_T_1 == 8'hFB & write_0_en];
      Register_inst252 <= _T_254[_T_1 == 8'hFC & write_0_en];
      Register_inst253 <= _T_255[_T_1 == 8'hFD & write_0_en];
      Register_inst254 <= _T_256[_T_1 == 8'hFE & write_0_en];
      Register_inst255 <= _T_257[&_T_1 & write_0_en];
    end
  end // always_ff @(posedge or posedge)
  initial begin
    Register_inst0 = 32'h0;
    Register_inst1 = 32'h0;
    Register_inst2 = 32'h0;
    Register_inst3 = 32'h0;
    Register_inst4 = 32'h0;
    Register_inst5 = 32'h0;
    Register_inst6 = 32'h0;
    Register_inst7 = 32'h0;
    Register_inst8 = 32'h0;
    Register_inst9 = 32'h0;
    Register_inst10 = 32'h0;
    Register_inst11 = 32'h0;
    Register_inst12 = 32'h0;
    Register_inst13 = 32'h0;
    Register_inst14 = 32'h0;
    Register_inst15 = 32'h0;
    Register_inst16 = 32'h0;
    Register_inst17 = 32'h0;
    Register_inst18 = 32'h0;
    Register_inst19 = 32'h0;
    Register_inst20 = 32'h0;
    Register_inst21 = 32'h0;
    Register_inst22 = 32'h0;
    Register_inst23 = 32'h0;
    Register_inst24 = 32'h0;
    Register_inst25 = 32'h0;
    Register_inst26 = 32'h0;
    Register_inst27 = 32'h0;
    Register_inst28 = 32'h0;
    Register_inst29 = 32'h0;
    Register_inst30 = 32'h0;
    Register_inst31 = 32'h0;
    Register_inst32 = 32'h0;
    Register_inst33 = 32'h0;
    Register_inst34 = 32'h0;
    Register_inst35 = 32'h0;
    Register_inst36 = 32'h0;
    Register_inst37 = 32'h0;
    Register_inst38 = 32'h0;
    Register_inst39 = 32'h0;
    Register_inst40 = 32'h0;
    Register_inst41 = 32'h0;
    Register_inst42 = 32'h0;
    Register_inst43 = 32'h0;
    Register_inst44 = 32'h0;
    Register_inst45 = 32'h0;
    Register_inst46 = 32'h0;
    Register_inst47 = 32'h0;
    Register_inst48 = 32'h0;
    Register_inst49 = 32'h0;
    Register_inst50 = 32'h0;
    Register_inst51 = 32'h0;
    Register_inst52 = 32'h0;
    Register_inst53 = 32'h0;
    Register_inst54 = 32'h0;
    Register_inst55 = 32'h0;
    Register_inst56 = 32'h0;
    Register_inst57 = 32'h0;
    Register_inst58 = 32'h0;
    Register_inst59 = 32'h0;
    Register_inst60 = 32'h0;
    Register_inst61 = 32'h0;
    Register_inst62 = 32'h0;
    Register_inst63 = 32'h0;
    Register_inst64 = 32'h0;
    Register_inst65 = 32'h0;
    Register_inst66 = 32'h0;
    Register_inst67 = 32'h0;
    Register_inst68 = 32'h0;
    Register_inst69 = 32'h0;
    Register_inst70 = 32'h0;
    Register_inst71 = 32'h0;
    Register_inst72 = 32'h0;
    Register_inst73 = 32'h0;
    Register_inst74 = 32'h0;
    Register_inst75 = 32'h0;
    Register_inst76 = 32'h0;
    Register_inst77 = 32'h0;
    Register_inst78 = 32'h0;
    Register_inst79 = 32'h0;
    Register_inst80 = 32'h0;
    Register_inst81 = 32'h0;
    Register_inst82 = 32'h0;
    Register_inst83 = 32'h0;
    Register_inst84 = 32'h0;
    Register_inst85 = 32'h0;
    Register_inst86 = 32'h0;
    Register_inst87 = 32'h0;
    Register_inst88 = 32'h0;
    Register_inst89 = 32'h0;
    Register_inst90 = 32'h0;
    Register_inst91 = 32'h0;
    Register_inst92 = 32'h0;
    Register_inst93 = 32'h0;
    Register_inst94 = 32'h0;
    Register_inst95 = 32'h0;
    Register_inst96 = 32'h0;
    Register_inst97 = 32'h0;
    Register_inst98 = 32'h0;
    Register_inst99 = 32'h0;
    Register_inst100 = 32'h0;
    Register_inst101 = 32'h0;
    Register_inst102 = 32'h0;
    Register_inst103 = 32'h0;
    Register_inst104 = 32'h0;
    Register_inst105 = 32'h0;
    Register_inst106 = 32'h0;
    Register_inst107 = 32'h0;
    Register_inst108 = 32'h0;
    Register_inst109 = 32'h0;
    Register_inst110 = 32'h0;
    Register_inst111 = 32'h0;
    Register_inst112 = 32'h0;
    Register_inst113 = 32'h0;
    Register_inst114 = 32'h0;
    Register_inst115 = 32'h0;
    Register_inst116 = 32'h0;
    Register_inst117 = 32'h0;
    Register_inst118 = 32'h0;
    Register_inst119 = 32'h0;
    Register_inst120 = 32'h0;
    Register_inst121 = 32'h0;
    Register_inst122 = 32'h0;
    Register_inst123 = 32'h0;
    Register_inst124 = 32'h0;
    Register_inst125 = 32'h0;
    Register_inst126 = 32'h0;
    Register_inst127 = 32'h0;
    Register_inst128 = 32'h0;
    Register_inst129 = 32'h0;
    Register_inst130 = 32'h0;
    Register_inst131 = 32'h0;
    Register_inst132 = 32'h0;
    Register_inst133 = 32'h0;
    Register_inst134 = 32'h0;
    Register_inst135 = 32'h0;
    Register_inst136 = 32'h0;
    Register_inst137 = 32'h0;
    Register_inst138 = 32'h0;
    Register_inst139 = 32'h0;
    Register_inst140 = 32'h0;
    Register_inst141 = 32'h0;
    Register_inst142 = 32'h0;
    Register_inst143 = 32'h0;
    Register_inst144 = 32'h0;
    Register_inst145 = 32'h0;
    Register_inst146 = 32'h0;
    Register_inst147 = 32'h0;
    Register_inst148 = 32'h0;
    Register_inst149 = 32'h0;
    Register_inst150 = 32'h0;
    Register_inst151 = 32'h0;
    Register_inst152 = 32'h0;
    Register_inst153 = 32'h0;
    Register_inst154 = 32'h0;
    Register_inst155 = 32'h0;
    Register_inst156 = 32'h0;
    Register_inst157 = 32'h0;
    Register_inst158 = 32'h0;
    Register_inst159 = 32'h0;
    Register_inst160 = 32'h0;
    Register_inst161 = 32'h0;
    Register_inst162 = 32'h0;
    Register_inst163 = 32'h0;
    Register_inst164 = 32'h0;
    Register_inst165 = 32'h0;
    Register_inst166 = 32'h0;
    Register_inst167 = 32'h0;
    Register_inst168 = 32'h0;
    Register_inst169 = 32'h0;
    Register_inst170 = 32'h0;
    Register_inst171 = 32'h0;
    Register_inst172 = 32'h0;
    Register_inst173 = 32'h0;
    Register_inst174 = 32'h0;
    Register_inst175 = 32'h0;
    Register_inst176 = 32'h0;
    Register_inst177 = 32'h0;
    Register_inst178 = 32'h0;
    Register_inst179 = 32'h0;
    Register_inst180 = 32'h0;
    Register_inst181 = 32'h0;
    Register_inst182 = 32'h0;
    Register_inst183 = 32'h0;
    Register_inst184 = 32'h0;
    Register_inst185 = 32'h0;
    Register_inst186 = 32'h0;
    Register_inst187 = 32'h0;
    Register_inst188 = 32'h0;
    Register_inst189 = 32'h0;
    Register_inst190 = 32'h0;
    Register_inst191 = 32'h0;
    Register_inst192 = 32'h0;
    Register_inst193 = 32'h0;
    Register_inst194 = 32'h0;
    Register_inst195 = 32'h0;
    Register_inst196 = 32'h0;
    Register_inst197 = 32'h0;
    Register_inst198 = 32'h0;
    Register_inst199 = 32'h0;
    Register_inst200 = 32'h0;
    Register_inst201 = 32'h0;
    Register_inst202 = 32'h0;
    Register_inst203 = 32'h0;
    Register_inst204 = 32'h0;
    Register_inst205 = 32'h0;
    Register_inst206 = 32'h0;
    Register_inst207 = 32'h0;
    Register_inst208 = 32'h0;
    Register_inst209 = 32'h0;
    Register_inst210 = 32'h0;
    Register_inst211 = 32'h0;
    Register_inst212 = 32'h0;
    Register_inst213 = 32'h0;
    Register_inst214 = 32'h0;
    Register_inst215 = 32'h0;
    Register_inst216 = 32'h0;
    Register_inst217 = 32'h0;
    Register_inst218 = 32'h0;
    Register_inst219 = 32'h0;
    Register_inst220 = 32'h0;
    Register_inst221 = 32'h0;
    Register_inst222 = 32'h0;
    Register_inst223 = 32'h0;
    Register_inst224 = 32'h0;
    Register_inst225 = 32'h0;
    Register_inst226 = 32'h0;
    Register_inst227 = 32'h0;
    Register_inst228 = 32'h0;
    Register_inst229 = 32'h0;
    Register_inst230 = 32'h0;
    Register_inst231 = 32'h0;
    Register_inst232 = 32'h0;
    Register_inst233 = 32'h0;
    Register_inst234 = 32'h0;
    Register_inst235 = 32'h0;
    Register_inst236 = 32'h0;
    Register_inst237 = 32'h0;
    Register_inst238 = 32'h0;
    Register_inst239 = 32'h0;
    Register_inst240 = 32'h0;
    Register_inst241 = 32'h0;
    Register_inst242 = 32'h0;
    Register_inst243 = 32'h0;
    Register_inst244 = 32'h0;
    Register_inst245 = 32'h0;
    Register_inst246 = 32'h0;
    Register_inst247 = 32'h0;
    Register_inst248 = 32'h0;
    Register_inst249 = 32'h0;
    Register_inst250 = 32'h0;
    Register_inst251 = 32'h0;
    Register_inst252 = 32'h0;
    Register_inst253 = 32'h0;
    Register_inst254 = 32'h0;
    Register_inst255 = 32'h0;
  end // initial
  wire [255:0][31:0] _T = {{Register_inst0}, {Register_inst1}, {Register_inst2}, {Register_inst3}, {Register_inst4},
                {Register_inst5}, {Register_inst6}, {Register_inst7}, {Register_inst8}, {Register_inst9},
                {Register_inst10}, {Register_inst11}, {Register_inst12}, {Register_inst13},
                {Register_inst14}, {Register_inst15}, {Register_inst16}, {Register_inst17},
                {Register_inst18}, {Register_inst19}, {Register_inst20}, {Register_inst21},
                {Register_inst22}, {Register_inst23}, {Register_inst24}, {Register_inst25},
                {Register_inst26}, {Register_inst27}, {Register_inst28}, {Register_inst29},
                {Register_inst30}, {Register_inst31}, {Register_inst32}, {Register_inst33},
                {Register_inst34}, {Register_inst35}, {Register_inst36}, {Register_inst37},
                {Register_inst38}, {Register_inst39}, {Register_inst40}, {Register_inst41},
                {Register_inst42}, {Register_inst43}, {Register_inst44}, {Register_inst45},
                {Register_inst46}, {Register_inst47}, {Register_inst48}, {Register_inst49},
                {Register_inst50}, {Register_inst51}, {Register_inst52}, {Register_inst53},
                {Register_inst54}, {Register_inst55}, {Register_inst56}, {Register_inst57},
                {Register_inst58}, {Register_inst59}, {Register_inst60}, {Register_inst61},
                {Register_inst62}, {Register_inst63}, {Register_inst64}, {Register_inst65},
                {Register_inst66}, {Register_inst67}, {Register_inst68}, {Register_inst69},
                {Register_inst70}, {Register_inst71}, {Register_inst72}, {Register_inst73},
                {Register_inst74}, {Register_inst75}, {Register_inst76}, {Register_inst77},
                {Register_inst78}, {Register_inst79}, {Register_inst80}, {Register_inst81},
                {Register_inst82}, {Register_inst83}, {Register_inst84}, {Register_inst85},
                {Register_inst86}, {Register_inst87}, {Register_inst88}, {Register_inst89},
                {Register_inst90}, {Register_inst91}, {Register_inst92}, {Register_inst93},
                {Register_inst94}, {Register_inst95}, {Register_inst96}, {Register_inst97},
                {Register_inst98}, {Register_inst99}, {Register_inst100}, {Register_inst101},
                {Register_inst102}, {Register_inst103}, {Register_inst104}, {Register_inst105},
                {Register_inst106}, {Register_inst107}, {Register_inst108}, {Register_inst109},
                {Register_inst110}, {Register_inst111}, {Register_inst112}, {Register_inst113},
                {Register_inst114}, {Register_inst115}, {Register_inst116}, {Register_inst117},
                {Register_inst118}, {Register_inst119}, {Register_inst120}, {Register_inst121},
                {Register_inst122}, {Register_inst123}, {Register_inst124}, {Register_inst125},
                {Register_inst126}, {Register_inst127}, {Register_inst128}, {Register_inst129},
                {Register_inst130}, {Register_inst131}, {Register_inst132}, {Register_inst133},
                {Register_inst134}, {Register_inst135}, {Register_inst136}, {Register_inst137},
                {Register_inst138}, {Register_inst139}, {Register_inst140}, {Register_inst141},
                {Register_inst142}, {Register_inst143}, {Register_inst144}, {Register_inst145},
                {Register_inst146}, {Register_inst147}, {Register_inst148}, {Register_inst149},
                {Register_inst150}, {Register_inst151}, {Register_inst152}, {Register_inst153},
                {Register_inst154}, {Register_inst155}, {Register_inst156}, {Register_inst157},
                {Register_inst158}, {Register_inst159}, {Register_inst160}, {Register_inst161},
                {Register_inst162}, {Register_inst163}, {Register_inst164}, {Register_inst165},
                {Register_inst166}, {Register_inst167}, {Register_inst168}, {Register_inst169},
                {Register_inst170}, {Register_inst171}, {Register_inst172}, {Register_inst173},
                {Register_inst174}, {Register_inst175}, {Register_inst176}, {Register_inst177},
                {Register_inst178}, {Register_inst179}, {Register_inst180}, {Register_inst181},
                {Register_inst182}, {Register_inst183}, {Register_inst184}, {Register_inst185},
                {Register_inst186}, {Register_inst187}, {Register_inst188}, {Register_inst189},
                {Register_inst190}, {Register_inst191}, {Register_inst192}, {Register_inst193},
                {Register_inst194}, {Register_inst195}, {Register_inst196}, {Register_inst197},
                {Register_inst198}, {Register_inst199}, {Register_inst200}, {Register_inst201},
                {Register_inst202}, {Register_inst203}, {Register_inst204}, {Register_inst205},
                {Register_inst206}, {Register_inst207}, {Register_inst208}, {Register_inst209},
                {Register_inst210}, {Register_inst211}, {Register_inst212}, {Register_inst213},
                {Register_inst214}, {Register_inst215}, {Register_inst216}, {Register_inst217},
                {Register_inst218}, {Register_inst219}, {Register_inst220}, {Register_inst221},
                {Register_inst222}, {Register_inst223}, {Register_inst224}, {Register_inst225},
                {Register_inst226}, {Register_inst227}, {Register_inst228}, {Register_inst229},
                {Register_inst230}, {Register_inst231}, {Register_inst232}, {Register_inst233},
                {Register_inst234}, {Register_inst235}, {Register_inst236}, {Register_inst237},
                {Register_inst238}, {Register_inst239}, {Register_inst240}, {Register_inst241},
                {Register_inst242}, {Register_inst243}, {Register_inst244}, {Register_inst245},
                {Register_inst246}, {Register_inst247}, {Register_inst248}, {Register_inst249},
                {Register_inst250}, {Register_inst251}, {Register_inst252}, {Register_inst253},
                {Register_inst254}, {Register_inst255}};
  assign code_read_0_data = _T[code_read_0_addr];
endmodule

module Risc(
  input         is_write,
  input  [7:0]  write_addr,
  input  [31:0] write_data,
  input         boot, CLK, ASYNCRESET,
  output        valid,
  output [31:0] out);

  wire [31:0] _T;
  wire [31:0] file_file_read_0_data;
  wire [31:0] file_file_read_1_data;
  wire [31:0] code_code_read_0_data;
  reg  [7:0]  Register_inst0;

  always_ff @(posedge CLK) begin
    automatic logic [1:0][7:0] _T_11 = {{Register_inst0 + 8'h1}, {8'h0}};
    automatic logic [1:0][7:0] _T_12 = {{_T_11[boot]}, {Register_inst0}};

    Register_inst0 <= _T_12[is_write];
  end // always_ff @(posedge)
  initial
    Register_inst0 = 8'h0;
  wire struct packed {logic [31:0] data; logic [7:0] addr; } _T_0 = '{data: write_data, addr: write_addr};
  wire [1:0] _T_1 = {{1'h0}, {1'h1}};
  wire [1:0] _T_2 = {{_T_1[&(code_code_read_0_data[23:16])]}, {1'h0}};
  wire [1:0] _T_3 = {{_T_2[boot]}, {1'h0}};
  wire [1:0][31:0] _T_4 = {{32'h0}, {{24'h0, code_code_read_0_data[7:0]}}};
  wire struct packed {logic [31:0] data; logic [7:0] addr; } _T_5 = '{data: _T, addr: (code_code_read_0_data[23:16])};
  wire [1:0][31:0] _T_6 = {{file_file_read_0_data}, {32'h0}};
  wire [1:0][31:0] _T_7 = {{file_file_read_1_data}, {32'h0}};
  wire [1:0][31:0] _T_8 = {{_T_4[code_code_read_0_data[31:24] == 8'h1]}, {_T_6[code_code_read_0_data[15:8] == 8'h0] +
                _T_7[code_code_read_0_data[7:0] == 8'h0]}};
  wire [1:0][31:0] _T_9 = {{_T_8[code_code_read_0_data[31:24] == 8'h0]}, {32'h0}};
  wire [1:0][31:0] _T_10 = {{_T_9[boot]}, {32'h0}};
  assign _T = _T_10[is_write];
  code code (
    .CLK              (CLK),
    .ASYNCRESET       (ASYNCRESET),
    .code_read_0_addr (Register_inst0),
    .write_0          (_T_0),
    .write_0_en       (is_write),
    .code_read_0_data (code_code_read_0_data)
  );
  file file (
    .CLK              (CLK),
    .ASYNCRESET       (ASYNCRESET),
    .file_read_0_addr (code_code_read_0_data[15:8]),
    .file_read_1_addr (code_code_read_0_data[7:0]),
    .write_0          (_T_5),
    .write_0_en       (code_code_read_0_data[23:16] != 8'hFF),
    .file_read_0_data (file_file_read_0_data),
    .file_read_1_data (file_file_read_1_data)
  );
  assign valid = _T_3[is_write];
  assign out = _T;
endmodule

