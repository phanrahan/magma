module simple_comb(
  input  [15:0] a,
                b,
                c,
  output [15:0] y,
                z
);

  assign y = 16'hFFFF;
  assign z = 16'hFFFF;
endmodule

