module main (
    input [1:0] I,
    output [1:0] O
);
assign O = I;
endmodule

