module no_outputs(
  input I
);

endmodule

