module simple_mixed_direction_ports(	// <stdin>:1:1
  input  [7:0] a_x,
  output [7:0] a_y);

  assign a_y = a_x;	// <stdin>:2:5
endmodule

