module LUT(
  input  [7:0] I,
  output [7:0] O);

wire [255:0] _T = {{1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0},
                {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1},
                {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0},
                {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1},
                {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0},
                {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1},
                {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0},
                {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1},
                {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0},
                {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1},
                {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0},
                {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1},
                {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0},
                {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1},
                {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0},
                {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1},
                {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0},
                {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1},
                {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0},
                {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1},
                {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0},
                {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1},
                {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0}, {1'h1}, {1'h0},
                {1'h1}, {1'h0}, {1'h1}};
wire [255:0] _T_0 = {{1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1},
                {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0},
                {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0},
                {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1},
                {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1},
                {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0},
                {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0},
                {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1},
                {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1},
                {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0},
                {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0},
                {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1},
                {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1},
                {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0},
                {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0},
                {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1},
                {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1},
                {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0},
                {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0},
                {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1},
                {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1},
                {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0},
                {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h0},
                {1'h0}, {1'h1}, {1'h1}};
wire [255:0] _T_1 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}};
wire [255:0] _T_2 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}};
wire [255:0] _T_3 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}};
wire [255:0] _T_4 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}};
wire [255:0] _T_5 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}};
wire [255:0] _T_6 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0},
                {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1}, {1'h1},
                {1'h1}, {1'h1}, {1'h1}};
  assign O = {_T_6[I], _T_5[I], _T_4[I], _T_3[I], _T_2[I], _T_1[I], _T_0[I], _T[I]};
endmodule

module Tbl(
  input  [7:0] addr,
  output [7:0] out);

  LUT LUT_inst0 (
    .I (addr),
    .O (out)
  );
endmodule

