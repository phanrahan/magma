module LUT(
  input  [1:0] I,
  output [7:0] O);

  assign O = {({{1'h1}, {1'h1}, {1'h1}, {1'h1}})[I], ({{1'h1}, {1'h0}, {1'h0}, {1'h1}})[I], ({{1'h0}, {1'h1}, {1'h1}, {1'h1}})[I], ({{1'h1}, {1'h0}, {1'h1}, {1'h0}})[I], ({{1'h1}, {1'h1}, {1'h1}, {1'h1}})[I], ({{1'h1}, {1'h1}, {1'h1}, {1'h1}})[I], ({{1'h1}, {1'h0}, {1'h1}, {1'h1}})[I], ({{1'h0}, {1'h1}, {1'h0}, {1'h1}})[I]};	// <stdin>:3:13, :4:14, :5:10, :6:10, :7:10, :8:10, :9:10, :10:10, :11:10, :12:10, :13:10, :14:10, :15:11, :16:11, :17:11, :18:11, :19:11, :20:11, :21:11, :22:5
endmodule

module simple_lut(
  input  [1:0] a,
  output [7:0] y);

  LUT LUT_inst0 (	// <stdin>:25:20
    .I (a),
    .O (y)
  );
endmodule

