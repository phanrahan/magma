module simple_undriven(	// <stdin>:1:1
  output O);

  assign O = 1'bx;	// <stdin>:2:10, :4:5
endmodule

