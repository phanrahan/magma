module coreir_term #(
    parameter width = 1
) (
    input [width-1:0] in
);

endmodule

module MonitorWrapper (
    input [7:0] arr [63:0]
);
wire [7:0] MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0 [63:0];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[63] = arr[63];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[62] = arr[62];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[61] = arr[61];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[60] = arr[60];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[59] = arr[59];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[58] = arr[58];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[57] = arr[57];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[56] = arr[56];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[55] = arr[55];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[54] = arr[54];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[53] = arr[53];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[52] = arr[52];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[51] = arr[51];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[50] = arr[50];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[49] = arr[49];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[48] = arr[48];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[47] = arr[47];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[46] = arr[46];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[45] = arr[45];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[44] = arr[44];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[43] = arr[43];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[42] = arr[42];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[41] = arr[41];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[40] = arr[40];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[39] = arr[39];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[38] = arr[38];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[37] = arr[37];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[36] = arr[36];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[35] = arr[35];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[34] = arr[34];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[33] = arr[33];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[32] = arr[32];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[31] = arr[31];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[30] = arr[30];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[29] = arr[29];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[28] = arr[28];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[27] = arr[27];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[26] = arr[26];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[25] = arr[25];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[24] = arr[24];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[23] = arr[23];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[22] = arr[22];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[21] = arr[21];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[20] = arr[20];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[19] = arr[19];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[18] = arr[18];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[17] = arr[17];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[16] = arr[16];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[15] = arr[15];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[14] = arr[14];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[13] = arr[13];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[12] = arr[12];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[11] = arr[11];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[10] = arr[10];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[9] = arr[9];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[8] = arr[8];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[7] = arr[7];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[6] = arr[6];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[5] = arr[5];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[4] = arr[4];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[3] = arr[3];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[2] = arr[2];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[1] = arr[1];
assign MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0[0] = arr[0];

monitor #(.WIDTH(8), .DEPTH(64)) monitor_inst(.arr(MonitorWrapper_inline_verilog_inst_0___magma_inline_value_0));
                    
endmodule

