module Top(
  input  I,
  output O
);

  wire _magma_bind_wire_0 = I;
  assign O = I;
endmodule

