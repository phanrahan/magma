module mantle_sliceArrT__hi4__lo2__t_0BitIn_1BitIn24 (
    input in_0__0,
    input [1:0] in_0__1,
    input in_1__0,
    input [1:0] in_1__1,
    input in_2__0,
    input [1:0] in_2__1,
    input in_3__0,
    input [1:0] in_3__1,
    output out_0__0,
    output [1:0] out_0__1,
    output out_1__0,
    output [1:0] out_1__1
);
assign out_0__0 = in_2__0;
assign out_0__1 = in_2__1;
assign out_1__0 = in_3__0;
assign out_1__1 = in_3__1;
endmodule

module mantle_sliceArrT__hi2__lo0__t_0BitIn_1BitIn24 (
    input in_0__0,
    input [1:0] in_0__1,
    input in_1__0,
    input [1:0] in_1__1,
    input in_2__0,
    input [1:0] in_2__1,
    input in_3__0,
    input [1:0] in_3__1,
    output out_0__0,
    output [1:0] out_0__1,
    output out_1__0,
    output [1:0] out_1__1
);
assign out_0__0 = in_0__0;
assign out_0__1 = in_0__1;
assign out_1__0 = in_1__0;
assign out_1__1 = in_1__1;
endmodule

module mantle_liftArrT__t_0Bit_1Bit21 (
    input in__0,
    input [1:0] in__1,
    output out_0__0,
    output [1:0] out_0__1
);
assign out_0__0 = in__0;
assign out_0__1 = in__1;
endmodule

module mantle_getArrT__i3__t_0BitIn_1BitIn24 (
    input in_0__0,
    input [1:0] in_0__1,
    input in_1__0,
    input [1:0] in_1__1,
    input in_2__0,
    input [1:0] in_2__1,
    input in_3__0,
    input [1:0] in_3__1,
    output out__0,
    output [1:0] out__1
);
assign out__0 = in_3__0;
assign out__1 = in_3__1;
endmodule

module mantle_getArrT__i2__t_0BitIn_1BitIn24 (
    input in_0__0,
    input [1:0] in_0__1,
    input in_1__0,
    input [1:0] in_1__1,
    input in_2__0,
    input [1:0] in_2__1,
    input in_3__0,
    input [1:0] in_3__1,
    output out__0,
    output [1:0] out__1
);
assign out__0 = in_2__0;
assign out__1 = in_2__1;
endmodule

module mantle_getArrT__i1__t_0BitIn_1BitIn24 (
    input in_0__0,
    input [1:0] in_0__1,
    input in_1__0,
    input [1:0] in_1__1,
    input in_2__0,
    input [1:0] in_2__1,
    input in_3__0,
    input [1:0] in_3__1,
    output out__0,
    output [1:0] out__1
);
assign out__0 = in_1__0;
assign out__1 = in_1__1;
endmodule

module mantle_getArrT__i0__t_0BitIn_1BitIn24 (
    input in_0__0,
    input [1:0] in_0__1,
    input in_1__0,
    input [1:0] in_1__1,
    input in_2__0,
    input [1:0] in_2__1,
    input in_3__0,
    input [1:0] in_3__1,
    output out__0,
    output [1:0] out__1
);
assign out__0 = in_0__0;
assign out__1 = in_0__1;
endmodule

module mantle_concatArrT__t0_0BitIn_1BitIn22__t1_0BitIn_1BitIn22 (
    input in0_0__0,
    input [1:0] in0_0__1,
    input in0_1__0,
    input [1:0] in0_1__1,
    input in1_0__0,
    input [1:0] in1_0__1,
    input in1_1__0,
    input [1:0] in1_1__1,
    output out_0__0,
    output [1:0] out_0__1,
    output out_1__0,
    output [1:0] out_1__1,
    output out_2__0,
    output [1:0] out_2__1,
    output out_3__0,
    output [1:0] out_3__1
);
assign out_0__0 = in0_0__0;
assign out_0__1 = in0_0__1;
assign out_1__0 = in0_1__0;
assign out_1__1 = in0_1__1;
assign out_2__0 = in1_0__0;
assign out_2__1 = in1_0__1;
assign out_3__0 = in1_1__0;
assign out_3__1 = in1_1__1;
endmodule

module mantle_concatArrT__t0_0BitIn_1BitIn21__t1_0BitIn_1BitIn23 (
    input in0_0__0,
    input [1:0] in0_0__1,
    input in1_0__0,
    input [1:0] in1_0__1,
    input in1_1__0,
    input [1:0] in1_1__1,
    input in1_2__0,
    input [1:0] in1_2__1,
    output out_0__0,
    output [1:0] out_0__1,
    output out_1__0,
    output [1:0] out_1__1,
    output out_2__0,
    output [1:0] out_2__1,
    output out_3__0,
    output [1:0] out_3__1
);
assign out_0__0 = in0_0__0;
assign out_0__1 = in0_0__1;
assign out_1__0 = in1_0__0;
assign out_1__1 = in1_0__1;
assign out_2__0 = in1_1__0;
assign out_2__1 = in1_1__1;
assign out_3__0 = in1_2__0;
assign out_3__1 = in1_2__1;
endmodule

module mantle_concatArrT__t0_0BitIn_1BitIn21__t1_0BitIn_1BitIn22 (
    input in0_0__0,
    input [1:0] in0_0__1,
    input in1_0__0,
    input [1:0] in1_0__1,
    input in1_1__0,
    input [1:0] in1_1__1,
    output out_0__0,
    output [1:0] out_0__1,
    output out_1__0,
    output [1:0] out_1__1,
    output out_2__0,
    output [1:0] out_2__1
);
assign out_0__0 = in0_0__0;
assign out_0__1 = in0_0__1;
assign out_1__0 = in1_0__0;
assign out_1__1 = in1_0__1;
assign out_2__0 = in1_1__0;
assign out_2__1 = in1_1__1;
endmodule

module mantle_concatArrT__t0_0BitIn_1BitIn21__t1_0BitIn_1BitIn21 (
    input in0_0__0,
    input [1:0] in0_0__1,
    input in1_0__0,
    input [1:0] in1_0__1,
    output out_0__0,
    output [1:0] out_0__1,
    output out_1__0,
    output [1:0] out_1__1
);
assign out_0__0 = in0_0__0;
assign out_0__1 = in0_0__1;
assign out_1__0 = in1_0__0;
assign out_1__1 = in1_0__1;
endmodule

module Foo (
    input I_0__0,
    input [1:0] I_0__1,
    input I_1__0,
    input [1:0] I_1__1,
    input I_2__0,
    input [1:0] I_2__1,
    input I_3__0,
    input [1:0] I_3__1,
    output O0_0__0,
    output [1:0] O0_0__1,
    output O0_1__0,
    output [1:0] O0_1__1,
    output O0_2__0,
    output [1:0] O0_2__1,
    output O0_3__0,
    output [1:0] O0_3__1,
    output O1_0__0,
    output [1:0] O1_0__1,
    output O1_1__0,
    output [1:0] O1_1__1,
    output O1_2__0,
    output [1:0] O1_2__1,
    output O1_3__0,
    output [1:0] O1_3__1,
    output O2_0__0,
    output [1:0] O2_0__1,
    output O2_1__0,
    output [1:0] O2_1__1,
    output O2_2__0,
    output [1:0] O2_2__1,
    output O2_3__0,
    output [1:0] O2_3__1,
    output O3_0__0,
    output [1:0] O3_0__1,
    output O3_1__0,
    output [1:0] O3_1__1,
    output O3_2__0,
    output [1:0] O3_2__1,
    output O3_3__0,
    output [1:0] O3_3__1
);
wire Concat_inst0_out_0__0;
wire [1:0] Concat_inst0_out_0__1;
wire Concat_inst0_out_1__0;
wire [1:0] Concat_inst0_out_1__1;
wire Concat_inst0_out_2__0;
wire [1:0] Concat_inst0_out_2__1;
wire Concat_inst0_out_3__0;
wire [1:0] Concat_inst0_out_3__1;
wire Concat_inst1_out_0__0;
wire [1:0] Concat_inst1_out_0__1;
wire Concat_inst1_out_1__0;
wire [1:0] Concat_inst1_out_1__1;
wire Concat_inst1_out_2__0;
wire [1:0] Concat_inst1_out_2__1;
wire Concat_inst1_out_3__0;
wire [1:0] Concat_inst1_out_3__1;
wire Concat_inst2_out_0__0;
wire [1:0] Concat_inst2_out_0__1;
wire Concat_inst2_out_1__0;
wire [1:0] Concat_inst2_out_1__1;
wire Concat_inst2_out_2__0;
wire [1:0] Concat_inst2_out_2__1;
wire Concat_inst3_out_0__0;
wire [1:0] Concat_inst3_out_0__1;
wire Concat_inst3_out_1__0;
wire [1:0] Concat_inst3_out_1__1;
wire Concat_inst4_out_0__0;
wire [1:0] Concat_inst4_out_0__1;
wire Concat_inst4_out_1__0;
wire [1:0] Concat_inst4_out_1__1;
wire Concat_inst4_out_2__0;
wire [1:0] Concat_inst4_out_2__1;
wire Concat_inst4_out_3__0;
wire [1:0] Concat_inst4_out_3__1;
wire Index_inst0_out__0;
wire [1:0] Index_inst0_out__1;
wire Index_inst1_out__0;
wire [1:0] Index_inst1_out__1;
wire Index_inst2_out__0;
wire [1:0] Index_inst2_out__1;
wire Index_inst3_out__0;
wire [1:0] Index_inst3_out__1;
wire Lift_inst0_out_0__0;
wire [1:0] Lift_inst0_out_0__1;
wire Lift_inst1_out_0__0;
wire [1:0] Lift_inst1_out_0__1;
wire Lift_inst2_out_0__0;
wire [1:0] Lift_inst2_out_0__1;
wire Lift_inst3_out_0__0;
wire [1:0] Lift_inst3_out_0__1;
wire Slice_inst0_out_0__0;
wire [1:0] Slice_inst0_out_0__1;
wire Slice_inst0_out_1__0;
wire [1:0] Slice_inst0_out_1__1;
wire Slice_inst1_out_0__0;
wire [1:0] Slice_inst1_out_0__1;
wire Slice_inst1_out_1__0;
wire [1:0] Slice_inst1_out_1__1;
wire Slice_inst2_out_0__0;
wire [1:0] Slice_inst2_out_0__1;
wire Slice_inst2_out_1__0;
wire [1:0] Slice_inst2_out_1__1;
wire Slice_inst3_out_0__0;
wire [1:0] Slice_inst3_out_0__1;
wire Slice_inst3_out_1__0;
wire [1:0] Slice_inst3_out_1__1;
mantle_concatArrT__t0_0BitIn_1BitIn22__t1_0BitIn_1BitIn22 Concat_inst0 (
    .in0_0__0(Slice_inst0_out_0__0),
    .in0_0__1(Slice_inst0_out_0__1),
    .in0_1__0(Slice_inst0_out_1__0),
    .in0_1__1(Slice_inst0_out_1__1),
    .in1_0__0(Slice_inst1_out_0__0),
    .in1_0__1(Slice_inst1_out_0__1),
    .in1_1__0(Slice_inst1_out_1__0),
    .in1_1__1(Slice_inst1_out_1__1),
    .out_0__0(Concat_inst0_out_0__0),
    .out_0__1(Concat_inst0_out_0__1),
    .out_1__0(Concat_inst0_out_1__0),
    .out_1__1(Concat_inst0_out_1__1),
    .out_2__0(Concat_inst0_out_2__0),
    .out_2__1(Concat_inst0_out_2__1),
    .out_3__0(Concat_inst0_out_3__0),
    .out_3__1(Concat_inst0_out_3__1)
);
mantle_concatArrT__t0_0BitIn_1BitIn21__t1_0BitIn_1BitIn23 Concat_inst1 (
    .in0_0__0(Lift_inst0_out_0__0),
    .in0_0__1(Lift_inst0_out_0__1),
    .in1_0__0(Concat_inst2_out_0__0),
    .in1_0__1(Concat_inst2_out_0__1),
    .in1_1__0(Concat_inst2_out_1__0),
    .in1_1__1(Concat_inst2_out_1__1),
    .in1_2__0(Concat_inst2_out_2__0),
    .in1_2__1(Concat_inst2_out_2__1),
    .out_0__0(Concat_inst1_out_0__0),
    .out_0__1(Concat_inst1_out_0__1),
    .out_1__0(Concat_inst1_out_1__0),
    .out_1__1(Concat_inst1_out_1__1),
    .out_2__0(Concat_inst1_out_2__0),
    .out_2__1(Concat_inst1_out_2__1),
    .out_3__0(Concat_inst1_out_3__0),
    .out_3__1(Concat_inst1_out_3__1)
);
mantle_concatArrT__t0_0BitIn_1BitIn21__t1_0BitIn_1BitIn22 Concat_inst2 (
    .in0_0__0(Lift_inst1_out_0__0),
    .in0_0__1(Lift_inst1_out_0__1),
    .in1_0__0(Concat_inst3_out_0__0),
    .in1_0__1(Concat_inst3_out_0__1),
    .in1_1__0(Concat_inst3_out_1__0),
    .in1_1__1(Concat_inst3_out_1__1),
    .out_0__0(Concat_inst2_out_0__0),
    .out_0__1(Concat_inst2_out_0__1),
    .out_1__0(Concat_inst2_out_1__0),
    .out_1__1(Concat_inst2_out_1__1),
    .out_2__0(Concat_inst2_out_2__0),
    .out_2__1(Concat_inst2_out_2__1)
);
mantle_concatArrT__t0_0BitIn_1BitIn21__t1_0BitIn_1BitIn21 Concat_inst3 (
    .in0_0__0(Lift_inst2_out_0__0),
    .in0_0__1(Lift_inst2_out_0__1),
    .in1_0__0(Lift_inst3_out_0__0),
    .in1_0__1(Lift_inst3_out_0__1),
    .out_0__0(Concat_inst3_out_0__0),
    .out_0__1(Concat_inst3_out_0__1),
    .out_1__0(Concat_inst3_out_1__0),
    .out_1__1(Concat_inst3_out_1__1)
);
mantle_concatArrT__t0_0BitIn_1BitIn22__t1_0BitIn_1BitIn22 Concat_inst4 (
    .in0_0__0(Slice_inst2_out_0__0),
    .in0_0__1(Slice_inst2_out_0__1),
    .in0_1__0(Slice_inst2_out_1__0),
    .in0_1__1(Slice_inst2_out_1__1),
    .in1_0__0(Slice_inst3_out_0__0),
    .in1_0__1(Slice_inst3_out_0__1),
    .in1_1__0(Slice_inst3_out_1__0),
    .in1_1__1(Slice_inst3_out_1__1),
    .out_0__0(Concat_inst4_out_0__0),
    .out_0__1(Concat_inst4_out_0__1),
    .out_1__0(Concat_inst4_out_1__0),
    .out_1__1(Concat_inst4_out_1__1),
    .out_2__0(Concat_inst4_out_2__0),
    .out_2__1(Concat_inst4_out_2__1),
    .out_3__0(Concat_inst4_out_3__0),
    .out_3__1(Concat_inst4_out_3__1)
);
mantle_getArrT__i1__t_0BitIn_1BitIn24 Index_inst0 (
    .in_0__0(I_0__0),
    .in_0__1(I_0__1),
    .in_1__0(I_1__0),
    .in_1__1(I_1__1),
    .in_2__0(I_2__0),
    .in_2__1(I_2__1),
    .in_3__0(I_3__0),
    .in_3__1(I_3__1),
    .out__0(Index_inst0_out__0),
    .out__1(Index_inst0_out__1)
);
mantle_getArrT__i0__t_0BitIn_1BitIn24 Index_inst1 (
    .in_0__0(I_0__0),
    .in_0__1(I_0__1),
    .in_1__0(I_1__0),
    .in_1__1(I_1__1),
    .in_2__0(I_2__0),
    .in_2__1(I_2__1),
    .in_3__0(I_3__0),
    .in_3__1(I_3__1),
    .out__0(Index_inst1_out__0),
    .out__1(Index_inst1_out__1)
);
mantle_getArrT__i3__t_0BitIn_1BitIn24 Index_inst2 (
    .in_0__0(I_0__0),
    .in_0__1(I_0__1),
    .in_1__0(I_1__0),
    .in_1__1(I_1__1),
    .in_2__0(I_2__0),
    .in_2__1(I_2__1),
    .in_3__0(I_3__0),
    .in_3__1(I_3__1),
    .out__0(Index_inst2_out__0),
    .out__1(Index_inst2_out__1)
);
mantle_getArrT__i2__t_0BitIn_1BitIn24 Index_inst3 (
    .in_0__0(I_0__0),
    .in_0__1(I_0__1),
    .in_1__0(I_1__0),
    .in_1__1(I_1__1),
    .in_2__0(I_2__0),
    .in_2__1(I_2__1),
    .in_3__0(I_3__0),
    .in_3__1(I_3__1),
    .out__0(Index_inst3_out__0),
    .out__1(Index_inst3_out__1)
);
mantle_liftArrT__t_0Bit_1Bit21 Lift_inst0 (
    .in__0(Index_inst0_out__0),
    .in__1(Index_inst0_out__1),
    .out_0__0(Lift_inst0_out_0__0),
    .out_0__1(Lift_inst0_out_0__1)
);
mantle_liftArrT__t_0Bit_1Bit21 Lift_inst1 (
    .in__0(Index_inst1_out__0),
    .in__1(Index_inst1_out__1),
    .out_0__0(Lift_inst1_out_0__0),
    .out_0__1(Lift_inst1_out_0__1)
);
mantle_liftArrT__t_0Bit_1Bit21 Lift_inst2 (
    .in__0(Index_inst2_out__0),
    .in__1(Index_inst2_out__1),
    .out_0__0(Lift_inst2_out_0__0),
    .out_0__1(Lift_inst2_out_0__1)
);
mantle_liftArrT__t_0Bit_1Bit21 Lift_inst3 (
    .in__0(Index_inst3_out__0),
    .in__1(Index_inst3_out__1),
    .out_0__0(Lift_inst3_out_0__0),
    .out_0__1(Lift_inst3_out_0__1)
);
mantle_sliceArrT__hi4__lo2__t_0BitIn_1BitIn24 Slice_inst0 (
    .in_0__0(I_0__0),
    .in_0__1(I_0__1),
    .in_1__0(I_1__0),
    .in_1__1(I_1__1),
    .in_2__0(I_2__0),
    .in_2__1(I_2__1),
    .in_3__0(I_3__0),
    .in_3__1(I_3__1),
    .out_0__0(Slice_inst0_out_0__0),
    .out_0__1(Slice_inst0_out_0__1),
    .out_1__0(Slice_inst0_out_1__0),
    .out_1__1(Slice_inst0_out_1__1)
);
mantle_sliceArrT__hi2__lo0__t_0BitIn_1BitIn24 Slice_inst1 (
    .in_0__0(I_0__0),
    .in_0__1(I_0__1),
    .in_1__0(I_1__0),
    .in_1__1(I_1__1),
    .in_2__0(I_2__0),
    .in_2__1(I_2__1),
    .in_3__0(I_3__0),
    .in_3__1(I_3__1),
    .out_0__0(Slice_inst1_out_0__0),
    .out_0__1(Slice_inst1_out_0__1),
    .out_1__0(Slice_inst1_out_1__0),
    .out_1__1(Slice_inst1_out_1__1)
);
mantle_sliceArrT__hi4__lo2__t_0BitIn_1BitIn24 Slice_inst2 (
    .in_0__0(I_0__0),
    .in_0__1(I_0__1),
    .in_1__0(I_1__0),
    .in_1__1(I_1__1),
    .in_2__0(I_2__0),
    .in_2__1(I_2__1),
    .in_3__0(I_3__0),
    .in_3__1(I_3__1),
    .out_0__0(Slice_inst2_out_0__0),
    .out_0__1(Slice_inst2_out_0__1),
    .out_1__0(Slice_inst2_out_1__0),
    .out_1__1(Slice_inst2_out_1__1)
);
mantle_sliceArrT__hi2__lo0__t_0BitIn_1BitIn24 Slice_inst3 (
    .in_0__0(I_0__0),
    .in_0__1(I_0__1),
    .in_1__0(I_1__0),
    .in_1__1(I_1__1),
    .in_2__0(I_2__0),
    .in_2__1(I_2__1),
    .in_3__0(I_3__0),
    .in_3__1(I_3__1),
    .out_0__0(Slice_inst3_out_0__0),
    .out_0__1(Slice_inst3_out_0__1),
    .out_1__0(Slice_inst3_out_1__0),
    .out_1__1(Slice_inst3_out_1__1)
);
assign O0_0__0 = I_0__0;
assign O0_0__1 = I_0__1;
assign O0_1__0 = I_1__0;
assign O0_1__1 = I_1__1;
assign O0_2__0 = I_2__0;
assign O0_2__1 = I_2__1;
assign O0_3__0 = I_3__0;
assign O0_3__1 = I_3__1;
assign O1_0__0 = Concat_inst0_out_0__0;
assign O1_0__1 = Concat_inst0_out_0__1;
assign O1_1__0 = Concat_inst0_out_1__0;
assign O1_1__1 = Concat_inst0_out_1__1;
assign O1_2__0 = Concat_inst0_out_2__0;
assign O1_2__1 = Concat_inst0_out_2__1;
assign O1_3__0 = Concat_inst0_out_3__0;
assign O1_3__1 = Concat_inst0_out_3__1;
assign O2_0__0 = Concat_inst1_out_0__0;
assign O2_0__1 = Concat_inst1_out_0__1;
assign O2_1__0 = Concat_inst1_out_1__0;
assign O2_1__1 = Concat_inst1_out_1__1;
assign O2_2__0 = Concat_inst1_out_2__0;
assign O2_2__1 = Concat_inst1_out_2__1;
assign O2_3__0 = Concat_inst1_out_3__0;
assign O2_3__1 = Concat_inst1_out_3__1;
assign O3_0__0 = Concat_inst4_out_0__0;
assign O3_0__1 = Concat_inst4_out_0__1;
assign O3_1__0 = Concat_inst4_out_1__0;
assign O3_1__1 = Concat_inst4_out_1__1;
assign O3_2__0 = Concat_inst4_out_2__0;
assign O3_2__1 = Concat_inst4_out_2__1;
assign O3_3__0 = Concat_inst4_out_3__0;
assign O3_3__1 = Concat_inst4_out_3__1;
endmodule

