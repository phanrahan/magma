module main (output [1:0] O);
assign O = 2'h2;
endmodule

