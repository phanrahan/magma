module mod2 #(parameter KRATOS_INSTANCE_ID = 24'sd23)
(
    input I
);

endmodule   // mod
