module simple_length_one_bits(
  input  I,
  output O
);

  assign O = I;
endmodule

