module CSRGen(
  input                                                   stall,
  input  [2:0]                                            cmd,
  input  [31:0]                                           I,
                                                          pc,
                                                          addr,
                                                          inst,
  input                                                   illegal,
  input  [1:0]                                            st_type,
  input  [2:0]                                            ld_type,
  input                                                   pc_check,
  input  struct packed {logic valid; logic [31:0] data; } host_fromhost,
  input                                                   CLK,
                                                          RESET,
  output [31:0]                                           O,
  output                                                  expt,
  output [31:0]                                           evec,
                                                          epc,
                                                          host_tohost
);

  wire [31:0]      _GEN;
  reg  [31:0]      Register_inst2;
  wire             not_stall = ~stall;
  wire             _GEN_0 = pc_check & addr[1];
  wire [1:0]       _GEN_1 = {{|(addr[1:0])}, {1'h0}};
  wire [1:0]       _GEN_2 = {{addr[0]}, {_GEN_1[ld_type == 3'h1]}};
  wire [1:0]       _GEN_3 = {{addr[0]}, {_GEN_2[ld_type == 3'h2]}};
  wire             _GEN_4 = _GEN_3[ld_type == 3'h4];
  wire [1:0]       _GEN_5 = {{|(addr[1:0])}, {1'h0}};
  wire [1:0]       _GEN_6 = {{addr[0]}, {_GEN_5[st_type == 2'h1]}};
  wire             _GEN_7 = _GEN_6[st_type == 2'h2];
  reg  [1:0]       Register_inst6;
  wire             _GEN_8 = inst[29:28] <= Register_inst6;
  wire             _GEN_9 = cmd == 3'h1 | cmd[1] & (|(inst[19:15]));
  wire             _GEN_10 = cmd == 3'h4;
  wire             _GEN_11 = _GEN_10 & ~(inst[20]) & ~(inst[28]);
  wire             _GEN_12 = _GEN_10 & inst[20] & ~(inst[28]);
  wire             _GEN_13 =
    illegal | _GEN_0 | _GEN_4 | _GEN_7 | (|(cmd[1:0]))
    & ({inst[31:20] == 12'h300,
        inst[31:20] == 12'h781,
        inst[31:20] == 12'h780,
        inst[31:20] == 12'h344,
        inst[31:20] == 12'h343,
        inst[31:20] == 12'h342,
        inst[31:20] == 12'h341,
        inst[31:20] == 12'h340,
        inst[31:20] == 12'h741,
        inst[31:20] == 12'h701,
        inst[31:20] == 12'h321,
        inst[31:20] == 12'h304,
        inst[31:20] == 12'h302,
        inst[31:20] == 12'h301,
        inst[31:20] == 12'hF10,
        inst[31:20] == 12'hF01,
        inst[31:20] == 12'hF00,
        inst[31:20] == 12'h982,
        inst[31:20] == 12'h981,
        inst[31:20] == 12'h980,
        inst[31:20] == 12'h902,
        inst[31:20] == 12'h901,
        inst[31:20] == 12'h900,
        inst[31:20] == 12'hC82,
        inst[31:20] == 12'hC81,
        inst[31:20] == 12'hC80,
        inst[31:20] == 12'hC02,
        inst[31:20] == 12'hC01,
        inst[31:20] == 12'hC00} == 29'h0 | ~_GEN_8) | _GEN_9
    & ((&(inst[31:30])) | inst[31:20] == 12'h301 | inst[31:20] == 12'h302) | _GEN_10
    & ~_GEN_8 | _GEN_11 | _GEN_12;
  reg  [31:0]      Register_inst16;
  reg  [31:0]      Register_inst17;
  reg              Register_inst8;
  reg  [1:0]       Register_inst7;
  reg              Register_inst9;
  wire             is_mbadaddr = _GEN_0 | _GEN_4 | _GEN_7;
  reg  [31:0]      Register_inst18;
  reg              Register_inst10;
  reg              Register_inst12;
  reg              Register_inst11;
  reg              Register_inst13;
  reg  [31:0]      Register_inst0;
  reg  [31:0]      Register_inst1;
  reg  [31:0]      _GEN_14;
  always_comb begin
    _GEN_14 = Register_inst1;
    if (&Register_inst0)
      _GEN_14 = Register_inst1 + 32'h1;
  end // always_comb
  reg  [31:0]      Register_inst14;
  reg  [31:0]      Register_inst15;
  reg  [31:0]      Register_inst19;
  reg  [31:0]      Register_inst20;
  reg  [31:0]      _GEN_15;
  always_comb begin
    _GEN_15 = Register_inst20;
    if (host_fromhost.valid)
      _GEN_15 = host_fromhost.data;
  end // always_comb
  wire             is_inst_ret = inst != 32'h13 & (~_GEN_13 | _GEN_11 | _GEN_12) & ~stall;
  reg  [31:0]      Register_inst4;
  reg  [31:0]      _GEN_16;
  always_comb begin
    _GEN_16 = Register_inst4;
    if (is_inst_ret)
      _GEN_16 = Register_inst4 + 32'h1;
  end // always_comb
  reg  [31:0]      Register_inst3;
  reg  [31:0]      _GEN_17;
  always_comb begin
    _GEN_17 = Register_inst3;
    if (&Register_inst2)
      _GEN_17 = Register_inst3 + 32'h1;
  end // always_comb
  wire             is_inst_reth = is_inst_ret & (&Register_inst4);
  reg  [31:0]      Register_inst5;
  reg  [31:0]      _GEN_18;
  always_comb begin
    _GEN_18 = Register_inst5;
    if (is_inst_reth)
      _GEN_18 = Register_inst5 + 32'h1;
  end // always_comb
  reg  [31:0]      _GEN_19;
  reg  [31:0]      _GEN_20;
  reg              _GEN_21;
  reg              _GEN_22;
  reg              _GEN_23;
  reg              _GEN_24;
  reg              _GEN_25;
  reg              _GEN_26;
  reg              _GEN_27;
  reg              _GEN_28;
  reg              _GEN_29;
  reg              _GEN_30;
  reg              _GEN_31;
  reg              _GEN_32;
  reg              _GEN_33;
  reg              _GEN_34;
  reg              _GEN_35;
  reg              _GEN_36;
  reg              _GEN_37;
  reg              _GEN_38;
  reg              _GEN_39;
  reg              _GEN_40;
  reg              _GEN_41;
  reg              _GEN_42;
  reg              _GEN_43;
  reg              _GEN_44;
  reg              _GEN_45;
  reg              _GEN_46;
  reg              _GEN_47;
  reg              _GEN_48;
  reg              _GEN_49;
  reg              _GEN_50;
  reg              _GEN_51;
  reg              _GEN_52;
  reg              _GEN_53;
  reg              _GEN_54;
  reg              _GEN_55;
  reg              _GEN_56;
  reg              _GEN_57;
  reg              _GEN_58;
  reg              _GEN_59;
  reg              _GEN_60;
  reg              _GEN_61;
  reg              _GEN_62;
  reg              _GEN_63;
  reg              _GEN_64;
  reg              _GEN_65;
  reg              _GEN_66;
  reg              _GEN_67;
  reg              _GEN_68;
  reg              _GEN_69;
  reg              _GEN_70;
  reg              _GEN_71;
  reg              _GEN_72;
  reg              _GEN_73;
  reg              _GEN_74;
  reg              _GEN_75;
  reg              _GEN_76;
  reg              _GEN_77;
  reg              _GEN_78;
  reg              _GEN_79;
  reg              _GEN_80;
  reg              _GEN_81;
  reg              _GEN_82;
  reg              _GEN_83;
  reg              _GEN_84;
  reg              _GEN_85;
  reg              _GEN_86;
  reg              _GEN_87;
  reg              _GEN_88;
  reg              _GEN_89;
  reg              _GEN_90;
  reg              _GEN_91;
  reg              _GEN_92;
  reg              _GEN_93;
  reg              _GEN_94;
  reg              _GEN_95;
  reg              _GEN_96;
  reg              _GEN_97;
  reg              _GEN_98;
  reg              _GEN_99;
  reg              _GEN_100;
  reg              _GEN_101;
  reg              _GEN_102;
  reg              _GEN_103;
  reg              _GEN_104;
  reg              _GEN_105;
  reg              _GEN_106;
  reg              _GEN_107;
  reg              _GEN_108;
  reg              _GEN_109;
  reg              _GEN_110;
  reg              _GEN_111;
  reg              _GEN_112;
  reg              _GEN_113;
  reg              _GEN_114;
  reg              _GEN_115;
  reg              _GEN_116;
  reg              _GEN_117;
  reg              _GEN_118;
  reg              _GEN_119;
  reg              _GEN_120;
  reg              _GEN_121;
  reg              _GEN_122;
  reg              _GEN_123;
  reg              _GEN_124;
  reg              _GEN_125;
  reg              _GEN_126;
  reg              _GEN_127;
  reg              _GEN_128;
  reg              _GEN_129;
  reg              _GEN_130;
  reg              _GEN_131;
  reg              _GEN_132;
  reg              _GEN_133;
  reg              _GEN_134;
  reg              _GEN_135;
  reg              _GEN_136;
  reg              _GEN_137;
  reg              _GEN_138;
  reg              _GEN_139;
  reg              _GEN_140;
  reg              _GEN_141;
  reg              _GEN_142;
  reg              _GEN_143;
  reg              _GEN_144;
  reg              _GEN_145;
  reg              _GEN_146;
  reg              _GEN_147;
  reg              _GEN_148;
  reg              _GEN_149;
  reg              _GEN_150;
  reg              _GEN_151;
  reg              _GEN_152;
  reg              _GEN_153;
  reg              _GEN_154;
  reg              _GEN_155;
  reg              _GEN_156;
  reg              _GEN_157;
  reg              _GEN_158;
  reg              _GEN_159;
  reg              _GEN_160;
  reg              _GEN_161;
  reg              _GEN_162;
  reg              _GEN_163;
  reg              _GEN_164;
  reg              _GEN_165;
  reg              _GEN_166;
  reg              _GEN_167;
  reg              _GEN_168;
  reg              _GEN_169;
  reg              _GEN_170;
  reg              _GEN_171;
  reg              _GEN_172;
  reg              _GEN_173;
  reg              _GEN_174;
  reg              _GEN_175;
  reg              _GEN_176;
  reg              _GEN_177;
  reg              _GEN_178;
  reg              _GEN_179;
  reg              _GEN_180;
  reg              _GEN_181;
  reg              _GEN_182;
  reg              _GEN_183;
  reg              _GEN_184;
  reg              _GEN_185;
  reg              _GEN_186;
  reg              _GEN_187;
  reg              _GEN_188;
  reg              _GEN_189;
  reg              _GEN_190;
  reg              _GEN_191;
  reg              _GEN_192;
  reg              _GEN_193;
  reg              _GEN_194;
  reg              _GEN_195;
  reg              _GEN_196;
  reg              _GEN_197;
  reg              _GEN_198;
  reg              _GEN_199;
  reg              _GEN_200;
  reg              _GEN_201;
  reg              _GEN_202;
  reg              _GEN_203;
  reg              _GEN_204;
  reg              _GEN_205;
  reg              _GEN_206;
  reg              _GEN_207;
  reg              _GEN_208;
  reg              _GEN_209;
  reg              _GEN_210;
  reg              _GEN_211;
  reg              _GEN_212;
  reg              _GEN_213;
  reg              _GEN_214;
  reg              _GEN_215;
  reg              _GEN_216;
  reg              _GEN_217;
  reg              _GEN_218;
  reg              _GEN_219;
  reg              _GEN_220;
  reg              _GEN_221;
  reg              _GEN_222;
  reg              _GEN_223;
  reg              _GEN_224;
  reg              _GEN_225;
  reg              _GEN_226;
  reg              _GEN_227;
  reg              _GEN_228;
  reg              _GEN_229;
  reg              _GEN_230;
  reg              _GEN_231;
  reg              _GEN_232;
  reg              _GEN_233;
  reg              _GEN_234;
  reg              _GEN_235;
  reg              _GEN_236;
  reg              _GEN_237;
  reg              _GEN_238;
  reg              _GEN_239;
  reg              _GEN_240;
  reg              _GEN_241;
  reg              _GEN_242;
  reg              _GEN_243;
  reg              _GEN_244;
  reg              _GEN_245;
  reg              _GEN_246;
  reg              _GEN_247;
  reg              _GEN_248;
  reg              _GEN_249;
  reg              _GEN_250;
  reg              _GEN_251;
  reg              _GEN_252;
  reg              _GEN_253;
  reg              _GEN_254;
  reg              _GEN_255;
  reg              _GEN_256;
  reg              _GEN_257;
  reg              _GEN_258;
  reg              _GEN_259;
  reg              _GEN_260;
  reg              _GEN_261;
  reg              _GEN_262;
  reg              _GEN_263;
  reg              _GEN_264;
  reg              _GEN_265;
  reg              _GEN_266;
  reg              _GEN_267;
  reg              _GEN_268;
  reg              _GEN_269;
  reg              _GEN_270;
  reg              _GEN_271;
  reg              _GEN_272;
  reg              _GEN_273;
  reg              _GEN_274;
  reg              _GEN_275;
  reg              _GEN_276;
  reg              _GEN_277;
  reg              _GEN_278;
  reg              _GEN_279;
  reg              _GEN_280;
  reg              _GEN_281;
  reg              _GEN_282;
  reg              _GEN_283;
  reg              _GEN_284;
  reg              _GEN_285;
  reg              _GEN_286;
  reg              _GEN_287;
  reg              _GEN_288;
  reg              _GEN_289;
  reg              _GEN_290;
  reg              _GEN_291;
  reg              _GEN_292;
  reg              _GEN_293;
  reg              _GEN_294;
  reg              _GEN_295;
  reg              _GEN_296;
  reg              _GEN_297;
  reg              _GEN_298;
  reg              _GEN_299;
  reg              _GEN_300;
  reg              _GEN_301;
  reg              _GEN_302;
  reg              _GEN_303;
  reg              _GEN_304;
  reg              _GEN_305;
  reg              _GEN_306;
  reg              _GEN_307;
  reg              _GEN_308;
  reg              _GEN_309;
  reg              _GEN_310;
  reg              _GEN_311;
  reg              _GEN_312;
  reg              _GEN_313;
  reg              _GEN_314;
  reg              _GEN_315;
  reg              _GEN_316;
  reg              _GEN_317;
  reg              _GEN_318;
  reg              _GEN_319;
  reg              _GEN_320;
  reg              _GEN_321;
  reg              _GEN_322;
  reg              _GEN_323;
  reg              _GEN_324;
  reg              _GEN_325;
  reg              _GEN_326;
  reg              _GEN_327;
  reg              _GEN_328;
  reg              _GEN_329;
  reg              _GEN_330;
  reg              _GEN_331;
  reg              _GEN_332;
  reg              _GEN_333;
  reg              _GEN_334;
  reg              _GEN_335;
  reg              _GEN_336;
  reg              _GEN_337;
  reg              _GEN_338;
  reg              _GEN_339;
  reg              _GEN_340;
  reg              _GEN_341;
  reg              _GEN_342;
  reg              _GEN_343;
  reg              _GEN_344;
  reg              _GEN_345;
  reg              _GEN_346;
  reg              _GEN_347;
  reg              _GEN_348;
  reg              _GEN_349;
  reg              _GEN_350;
  reg              _GEN_351;
  reg              _GEN_352;
  reg              _GEN_353;
  reg              _GEN_354;
  reg              _GEN_355;
  reg              _GEN_356;
  reg              _GEN_357;
  reg              _GEN_358;
  reg              _GEN_359;
  reg              _GEN_360;
  reg              _GEN_361;
  reg              _GEN_362;
  reg              _GEN_363;
  reg              _GEN_364;
  reg              _GEN_365;
  reg              _GEN_366;
  reg              _GEN_367;
  reg              _GEN_368;
  reg              _GEN_369;
  reg              _GEN_370;
  reg              _GEN_371;
  reg              _GEN_372;
  reg              _GEN_373;
  reg              _GEN_374;
  reg              _GEN_375;
  reg              _GEN_376;
  reg              _GEN_377;
  reg              _GEN_378;
  reg              _GEN_379;
  reg              _GEN_380;
  reg              _GEN_381;
  reg              _GEN_382;
  wire [1:0][31:0] _GEN_383 = {{I}, {32'h0}};
  wire [1:0][31:0] _GEN_384 = {{_GEN | I}, {_GEN_383[cmd == 3'h1]}};
  wire [1:0][31:0] _GEN_385 = {{_GEN & ~I}, {_GEN_384[cmd == 3'h2]}};
  wire [31:0]      _GEN_386 = _GEN_385[cmd == 3'h3];
  wire [31:0]      _GEN_387 = Register_inst0 + 32'h1;
  wire [31:0]      _GEN_388 = Register_inst2 + 32'h1;
  always_comb begin
    _GEN_19 = Register_inst16;
    _GEN_20 = Register_inst17;
    _GEN_21 = Register_inst6[0];
    _GEN_22 = Register_inst6[1];
    _GEN_23 = Register_inst8;
    _GEN_24 = Register_inst7[0];
    _GEN_25 = Register_inst7[1];
    _GEN_26 = Register_inst9;
    _GEN_27 = Register_inst18[0];
    _GEN_28 = Register_inst18[1];
    _GEN_29 = Register_inst18[2];
    _GEN_30 = Register_inst18[3];
    _GEN_31 = Register_inst18[4];
    _GEN_32 = Register_inst18[5];
    _GEN_33 = Register_inst18[6];
    _GEN_34 = Register_inst18[7];
    _GEN_35 = Register_inst18[8];
    _GEN_36 = Register_inst18[9];
    _GEN_37 = Register_inst18[10];
    _GEN_38 = Register_inst18[11];
    _GEN_39 = Register_inst18[12];
    _GEN_40 = Register_inst18[13];
    _GEN_41 = Register_inst18[14];
    _GEN_42 = Register_inst18[15];
    _GEN_43 = Register_inst18[16];
    _GEN_44 = Register_inst18[17];
    _GEN_45 = Register_inst18[18];
    _GEN_46 = Register_inst18[19];
    _GEN_47 = Register_inst18[20];
    _GEN_48 = Register_inst18[21];
    _GEN_49 = Register_inst18[22];
    _GEN_50 = Register_inst18[23];
    _GEN_51 = Register_inst18[24];
    _GEN_52 = Register_inst18[25];
    _GEN_53 = Register_inst18[26];
    _GEN_54 = Register_inst18[27];
    _GEN_55 = Register_inst18[28];
    _GEN_56 = Register_inst18[29];
    _GEN_57 = Register_inst18[30];
    _GEN_58 = Register_inst18[31];
    _GEN_59 = Register_inst10;
    _GEN_60 = Register_inst12;
    _GEN_61 = Register_inst11;
    _GEN_62 = Register_inst13;
    _GEN_63 = _GEN_387[0];
    _GEN_64 = _GEN_387[1];
    _GEN_65 = _GEN_387[2];
    _GEN_66 = _GEN_387[3];
    _GEN_67 = _GEN_387[4];
    _GEN_68 = _GEN_387[5];
    _GEN_69 = _GEN_387[6];
    _GEN_70 = _GEN_387[7];
    _GEN_71 = _GEN_387[8];
    _GEN_72 = _GEN_387[9];
    _GEN_73 = _GEN_387[10];
    _GEN_74 = _GEN_387[11];
    _GEN_75 = _GEN_387[12];
    _GEN_76 = _GEN_387[13];
    _GEN_77 = _GEN_387[14];
    _GEN_78 = _GEN_387[15];
    _GEN_79 = _GEN_387[16];
    _GEN_80 = _GEN_387[17];
    _GEN_81 = _GEN_387[18];
    _GEN_82 = _GEN_387[19];
    _GEN_83 = _GEN_387[20];
    _GEN_84 = _GEN_387[21];
    _GEN_85 = _GEN_387[22];
    _GEN_86 = _GEN_387[23];
    _GEN_87 = _GEN_387[24];
    _GEN_88 = _GEN_387[25];
    _GEN_89 = _GEN_387[26];
    _GEN_90 = _GEN_387[27];
    _GEN_91 = _GEN_387[28];
    _GEN_92 = _GEN_387[29];
    _GEN_93 = _GEN_387[30];
    _GEN_94 = _GEN_387[31];
    _GEN_95 = _GEN_14[0];
    _GEN_96 = _GEN_14[1];
    _GEN_97 = _GEN_14[2];
    _GEN_98 = _GEN_14[3];
    _GEN_99 = _GEN_14[4];
    _GEN_100 = _GEN_14[5];
    _GEN_101 = _GEN_14[6];
    _GEN_102 = _GEN_14[7];
    _GEN_103 = _GEN_14[8];
    _GEN_104 = _GEN_14[9];
    _GEN_105 = _GEN_14[10];
    _GEN_106 = _GEN_14[11];
    _GEN_107 = _GEN_14[12];
    _GEN_108 = _GEN_14[13];
    _GEN_109 = _GEN_14[14];
    _GEN_110 = _GEN_14[15];
    _GEN_111 = _GEN_14[16];
    _GEN_112 = _GEN_14[17];
    _GEN_113 = _GEN_14[18];
    _GEN_114 = _GEN_14[19];
    _GEN_115 = _GEN_14[20];
    _GEN_116 = _GEN_14[21];
    _GEN_117 = _GEN_14[22];
    _GEN_118 = _GEN_14[23];
    _GEN_119 = _GEN_14[24];
    _GEN_120 = _GEN_14[25];
    _GEN_121 = _GEN_14[26];
    _GEN_122 = _GEN_14[27];
    _GEN_123 = _GEN_14[28];
    _GEN_124 = _GEN_14[29];
    _GEN_125 = _GEN_14[30];
    _GEN_126 = _GEN_14[31];
    _GEN_127 = Register_inst14[0];
    _GEN_128 = Register_inst14[1];
    _GEN_129 = Register_inst14[2];
    _GEN_130 = Register_inst14[3];
    _GEN_131 = Register_inst14[4];
    _GEN_132 = Register_inst14[5];
    _GEN_133 = Register_inst14[6];
    _GEN_134 = Register_inst14[7];
    _GEN_135 = Register_inst14[8];
    _GEN_136 = Register_inst14[9];
    _GEN_137 = Register_inst14[10];
    _GEN_138 = Register_inst14[11];
    _GEN_139 = Register_inst14[12];
    _GEN_140 = Register_inst14[13];
    _GEN_141 = Register_inst14[14];
    _GEN_142 = Register_inst14[15];
    _GEN_143 = Register_inst14[16];
    _GEN_144 = Register_inst14[17];
    _GEN_145 = Register_inst14[18];
    _GEN_146 = Register_inst14[19];
    _GEN_147 = Register_inst14[20];
    _GEN_148 = Register_inst14[21];
    _GEN_149 = Register_inst14[22];
    _GEN_150 = Register_inst14[23];
    _GEN_151 = Register_inst14[24];
    _GEN_152 = Register_inst14[25];
    _GEN_153 = Register_inst14[26];
    _GEN_154 = Register_inst14[27];
    _GEN_155 = Register_inst14[28];
    _GEN_156 = Register_inst14[29];
    _GEN_157 = Register_inst14[30];
    _GEN_158 = Register_inst14[31];
    _GEN_159 = Register_inst15[0];
    _GEN_160 = Register_inst15[1];
    _GEN_161 = Register_inst15[2];
    _GEN_162 = Register_inst15[3];
    _GEN_163 = Register_inst15[4];
    _GEN_164 = Register_inst15[5];
    _GEN_165 = Register_inst15[6];
    _GEN_166 = Register_inst15[7];
    _GEN_167 = Register_inst15[8];
    _GEN_168 = Register_inst15[9];
    _GEN_169 = Register_inst15[10];
    _GEN_170 = Register_inst15[11];
    _GEN_171 = Register_inst15[12];
    _GEN_172 = Register_inst15[13];
    _GEN_173 = Register_inst15[14];
    _GEN_174 = Register_inst15[15];
    _GEN_175 = Register_inst15[16];
    _GEN_176 = Register_inst15[17];
    _GEN_177 = Register_inst15[18];
    _GEN_178 = Register_inst15[19];
    _GEN_179 = Register_inst15[20];
    _GEN_180 = Register_inst15[21];
    _GEN_181 = Register_inst15[22];
    _GEN_182 = Register_inst15[23];
    _GEN_183 = Register_inst15[24];
    _GEN_184 = Register_inst15[25];
    _GEN_185 = Register_inst15[26];
    _GEN_186 = Register_inst15[27];
    _GEN_187 = Register_inst15[28];
    _GEN_188 = Register_inst15[29];
    _GEN_189 = Register_inst15[30];
    _GEN_190 = Register_inst15[31];
    _GEN_191 = Register_inst19[0];
    _GEN_192 = Register_inst19[1];
    _GEN_193 = Register_inst19[2];
    _GEN_194 = Register_inst19[3];
    _GEN_195 = Register_inst19[4];
    _GEN_196 = Register_inst19[5];
    _GEN_197 = Register_inst19[6];
    _GEN_198 = Register_inst19[7];
    _GEN_199 = Register_inst19[8];
    _GEN_200 = Register_inst19[9];
    _GEN_201 = Register_inst19[10];
    _GEN_202 = Register_inst19[11];
    _GEN_203 = Register_inst19[12];
    _GEN_204 = Register_inst19[13];
    _GEN_205 = Register_inst19[14];
    _GEN_206 = Register_inst19[15];
    _GEN_207 = Register_inst19[16];
    _GEN_208 = Register_inst19[17];
    _GEN_209 = Register_inst19[18];
    _GEN_210 = Register_inst19[19];
    _GEN_211 = Register_inst19[20];
    _GEN_212 = Register_inst19[21];
    _GEN_213 = Register_inst19[22];
    _GEN_214 = Register_inst19[23];
    _GEN_215 = Register_inst19[24];
    _GEN_216 = Register_inst19[25];
    _GEN_217 = Register_inst19[26];
    _GEN_218 = Register_inst19[27];
    _GEN_219 = Register_inst19[28];
    _GEN_220 = Register_inst19[29];
    _GEN_221 = Register_inst19[30];
    _GEN_222 = Register_inst19[31];
    _GEN_223 = _GEN_15[0];
    _GEN_224 = _GEN_15[1];
    _GEN_225 = _GEN_15[2];
    _GEN_226 = _GEN_15[3];
    _GEN_227 = _GEN_15[4];
    _GEN_228 = _GEN_15[5];
    _GEN_229 = _GEN_15[6];
    _GEN_230 = _GEN_15[7];
    _GEN_231 = _GEN_15[8];
    _GEN_232 = _GEN_15[9];
    _GEN_233 = _GEN_15[10];
    _GEN_234 = _GEN_15[11];
    _GEN_235 = _GEN_15[12];
    _GEN_236 = _GEN_15[13];
    _GEN_237 = _GEN_15[14];
    _GEN_238 = _GEN_15[15];
    _GEN_239 = _GEN_15[16];
    _GEN_240 = _GEN_15[17];
    _GEN_241 = _GEN_15[18];
    _GEN_242 = _GEN_15[19];
    _GEN_243 = _GEN_15[20];
    _GEN_244 = _GEN_15[21];
    _GEN_245 = _GEN_15[22];
    _GEN_246 = _GEN_15[23];
    _GEN_247 = _GEN_15[24];
    _GEN_248 = _GEN_15[25];
    _GEN_249 = _GEN_15[26];
    _GEN_250 = _GEN_15[27];
    _GEN_251 = _GEN_15[28];
    _GEN_252 = _GEN_15[29];
    _GEN_253 = _GEN_15[30];
    _GEN_254 = _GEN_15[31];
    _GEN_255 = _GEN_388[0];
    _GEN_256 = _GEN_388[1];
    _GEN_257 = _GEN_388[2];
    _GEN_258 = _GEN_388[3];
    _GEN_259 = _GEN_388[4];
    _GEN_260 = _GEN_388[5];
    _GEN_261 = _GEN_388[6];
    _GEN_262 = _GEN_388[7];
    _GEN_263 = _GEN_388[8];
    _GEN_264 = _GEN_388[9];
    _GEN_265 = _GEN_388[10];
    _GEN_266 = _GEN_388[11];
    _GEN_267 = _GEN_388[12];
    _GEN_268 = _GEN_388[13];
    _GEN_269 = _GEN_388[14];
    _GEN_270 = _GEN_388[15];
    _GEN_271 = _GEN_388[16];
    _GEN_272 = _GEN_388[17];
    _GEN_273 = _GEN_388[18];
    _GEN_274 = _GEN_388[19];
    _GEN_275 = _GEN_388[20];
    _GEN_276 = _GEN_388[21];
    _GEN_277 = _GEN_388[22];
    _GEN_278 = _GEN_388[23];
    _GEN_279 = _GEN_388[24];
    _GEN_280 = _GEN_388[25];
    _GEN_281 = _GEN_388[26];
    _GEN_282 = _GEN_388[27];
    _GEN_283 = _GEN_388[28];
    _GEN_284 = _GEN_388[29];
    _GEN_285 = _GEN_388[30];
    _GEN_286 = _GEN_388[31];
    _GEN_287 = _GEN_16[0];
    _GEN_288 = _GEN_16[1];
    _GEN_289 = _GEN_16[2];
    _GEN_290 = _GEN_16[3];
    _GEN_291 = _GEN_16[4];
    _GEN_292 = _GEN_16[5];
    _GEN_293 = _GEN_16[6];
    _GEN_294 = _GEN_16[7];
    _GEN_295 = _GEN_16[8];
    _GEN_296 = _GEN_16[9];
    _GEN_297 = _GEN_16[10];
    _GEN_298 = _GEN_16[11];
    _GEN_299 = _GEN_16[12];
    _GEN_300 = _GEN_16[13];
    _GEN_301 = _GEN_16[14];
    _GEN_302 = _GEN_16[15];
    _GEN_303 = _GEN_16[16];
    _GEN_304 = _GEN_16[17];
    _GEN_305 = _GEN_16[18];
    _GEN_306 = _GEN_16[19];
    _GEN_307 = _GEN_16[20];
    _GEN_308 = _GEN_16[21];
    _GEN_309 = _GEN_16[22];
    _GEN_310 = _GEN_16[23];
    _GEN_311 = _GEN_16[24];
    _GEN_312 = _GEN_16[25];
    _GEN_313 = _GEN_16[26];
    _GEN_314 = _GEN_16[27];
    _GEN_315 = _GEN_16[28];
    _GEN_316 = _GEN_16[29];
    _GEN_317 = _GEN_16[30];
    _GEN_318 = _GEN_16[31];
    _GEN_319 = _GEN_17[0];
    _GEN_320 = _GEN_17[1];
    _GEN_321 = _GEN_17[2];
    _GEN_322 = _GEN_17[3];
    _GEN_323 = _GEN_17[4];
    _GEN_324 = _GEN_17[5];
    _GEN_325 = _GEN_17[6];
    _GEN_326 = _GEN_17[7];
    _GEN_327 = _GEN_17[8];
    _GEN_328 = _GEN_17[9];
    _GEN_329 = _GEN_17[10];
    _GEN_330 = _GEN_17[11];
    _GEN_331 = _GEN_17[12];
    _GEN_332 = _GEN_17[13];
    _GEN_333 = _GEN_17[14];
    _GEN_334 = _GEN_17[15];
    _GEN_335 = _GEN_17[16];
    _GEN_336 = _GEN_17[17];
    _GEN_337 = _GEN_17[18];
    _GEN_338 = _GEN_17[19];
    _GEN_339 = _GEN_17[20];
    _GEN_340 = _GEN_17[21];
    _GEN_341 = _GEN_17[22];
    _GEN_342 = _GEN_17[23];
    _GEN_343 = _GEN_17[24];
    _GEN_344 = _GEN_17[25];
    _GEN_345 = _GEN_17[26];
    _GEN_346 = _GEN_17[27];
    _GEN_347 = _GEN_17[28];
    _GEN_348 = _GEN_17[29];
    _GEN_349 = _GEN_17[30];
    _GEN_350 = _GEN_17[31];
    _GEN_351 = _GEN_18[0];
    _GEN_352 = _GEN_18[1];
    _GEN_353 = _GEN_18[2];
    _GEN_354 = _GEN_18[3];
    _GEN_355 = _GEN_18[4];
    _GEN_356 = _GEN_18[5];
    _GEN_357 = _GEN_18[6];
    _GEN_358 = _GEN_18[7];
    _GEN_359 = _GEN_18[8];
    _GEN_360 = _GEN_18[9];
    _GEN_361 = _GEN_18[10];
    _GEN_362 = _GEN_18[11];
    _GEN_363 = _GEN_18[12];
    _GEN_364 = _GEN_18[13];
    _GEN_365 = _GEN_18[14];
    _GEN_366 = _GEN_18[15];
    _GEN_367 = _GEN_18[16];
    _GEN_368 = _GEN_18[17];
    _GEN_369 = _GEN_18[18];
    _GEN_370 = _GEN_18[19];
    _GEN_371 = _GEN_18[20];
    _GEN_372 = _GEN_18[21];
    _GEN_373 = _GEN_18[22];
    _GEN_374 = _GEN_18[23];
    _GEN_375 = _GEN_18[24];
    _GEN_376 = _GEN_18[25];
    _GEN_377 = _GEN_18[26];
    _GEN_378 = _GEN_18[27];
    _GEN_379 = _GEN_18[28];
    _GEN_380 = _GEN_18[29];
    _GEN_381 = _GEN_18[30];
    _GEN_382 = _GEN_18[31];
    if (not_stall) begin
      if (_GEN_13) begin
        _GEN_19 = {pc[31:2], 2'h0};
        _GEN_21 = 1'h1;
        _GEN_22 = 1'h1;
        _GEN_23 = 1'h0;
        _GEN_24 = Register_inst6[0];
        _GEN_25 = Register_inst6[1];
        _GEN_26 = Register_inst8;
        if (_GEN_0)
          _GEN_20 = 32'h0;
        else if (_GEN_4)
          _GEN_20 = 32'h4;
        else if (_GEN_7)
          _GEN_20 = 32'h6;
        else if (_GEN_11)
          _GEN_20 = {30'h0, Register_inst6} + 32'h8;
        else if (_GEN_12)
          _GEN_20 = 32'h3;
        else
          _GEN_20 = 32'h2;
        if (is_mbadaddr) begin
          _GEN_27 = addr[0];
          _GEN_28 = addr[1];
          _GEN_29 = addr[2];
          _GEN_30 = addr[3];
          _GEN_31 = addr[4];
          _GEN_32 = addr[5];
          _GEN_33 = addr[6];
          _GEN_34 = addr[7];
          _GEN_35 = addr[8];
          _GEN_36 = addr[9];
          _GEN_37 = addr[10];
          _GEN_38 = addr[11];
          _GEN_39 = addr[12];
          _GEN_40 = addr[13];
          _GEN_41 = addr[14];
          _GEN_42 = addr[15];
          _GEN_43 = addr[16];
          _GEN_44 = addr[17];
          _GEN_45 = addr[18];
          _GEN_46 = addr[19];
          _GEN_47 = addr[20];
          _GEN_48 = addr[21];
          _GEN_49 = addr[22];
          _GEN_50 = addr[23];
          _GEN_51 = addr[24];
          _GEN_52 = addr[25];
          _GEN_53 = addr[26];
          _GEN_54 = addr[27];
          _GEN_55 = addr[28];
          _GEN_56 = addr[29];
          _GEN_57 = addr[30];
          _GEN_58 = addr[31];
        end
      end
      else if (_GEN_10 & ~(inst[20]) & inst[28]) begin
        _GEN_21 = Register_inst7[0];
        _GEN_22 = Register_inst7[1];
        _GEN_23 = Register_inst9;
        _GEN_24 = 1'h0;
        _GEN_25 = 1'h0;
        _GEN_26 = 1'h1;
      end
      else if (_GEN_9) begin
        if (inst[31:20] == 12'h300) begin
          _GEN_24 = _GEN_386[4];
          _GEN_25 = _GEN_386[5];
          _GEN_26 = _GEN_386[3];
          _GEN_21 = _GEN_386[1];
          _GEN_22 = _GEN_386[2];
          _GEN_23 = _GEN_386[0];
        end
        else if (inst[31:20] == 12'h344) begin
          _GEN_59 = _GEN_386[7];
          _GEN_60 = _GEN_386[3];
        end
        else if (inst[31:20] == 12'h304) begin
          _GEN_61 = _GEN_386[7];
          _GEN_62 = _GEN_386[3];
        end
        else if (inst[31:20] == 12'h701) begin
          _GEN_63 = _GEN_386[0];
          _GEN_64 = _GEN_386[1];
          _GEN_65 = _GEN_386[2];
          _GEN_66 = _GEN_386[3];
          _GEN_67 = _GEN_386[4];
          _GEN_68 = _GEN_386[5];
          _GEN_69 = _GEN_386[6];
          _GEN_70 = _GEN_386[7];
          _GEN_71 = _GEN_386[8];
          _GEN_72 = _GEN_386[9];
          _GEN_73 = _GEN_386[10];
          _GEN_74 = _GEN_386[11];
          _GEN_75 = _GEN_386[12];
          _GEN_76 = _GEN_386[13];
          _GEN_77 = _GEN_386[14];
          _GEN_78 = _GEN_386[15];
          _GEN_79 = _GEN_386[16];
          _GEN_80 = _GEN_386[17];
          _GEN_81 = _GEN_386[18];
          _GEN_82 = _GEN_386[19];
          _GEN_83 = _GEN_386[20];
          _GEN_84 = _GEN_386[21];
          _GEN_85 = _GEN_386[22];
          _GEN_86 = _GEN_386[23];
          _GEN_87 = _GEN_386[24];
          _GEN_88 = _GEN_386[25];
          _GEN_89 = _GEN_386[26];
          _GEN_90 = _GEN_386[27];
          _GEN_91 = _GEN_386[28];
          _GEN_92 = _GEN_386[29];
          _GEN_93 = _GEN_386[30];
          _GEN_94 = _GEN_386[31];
        end
        else if (inst[31:20] == 12'h741) begin
          _GEN_95 = _GEN_386[0];
          _GEN_96 = _GEN_386[1];
          _GEN_97 = _GEN_386[2];
          _GEN_98 = _GEN_386[3];
          _GEN_99 = _GEN_386[4];
          _GEN_100 = _GEN_386[5];
          _GEN_101 = _GEN_386[6];
          _GEN_102 = _GEN_386[7];
          _GEN_103 = _GEN_386[8];
          _GEN_104 = _GEN_386[9];
          _GEN_105 = _GEN_386[10];
          _GEN_106 = _GEN_386[11];
          _GEN_107 = _GEN_386[12];
          _GEN_108 = _GEN_386[13];
          _GEN_109 = _GEN_386[14];
          _GEN_110 = _GEN_386[15];
          _GEN_111 = _GEN_386[16];
          _GEN_112 = _GEN_386[17];
          _GEN_113 = _GEN_386[18];
          _GEN_114 = _GEN_386[19];
          _GEN_115 = _GEN_386[20];
          _GEN_116 = _GEN_386[21];
          _GEN_117 = _GEN_386[22];
          _GEN_118 = _GEN_386[23];
          _GEN_119 = _GEN_386[24];
          _GEN_120 = _GEN_386[25];
          _GEN_121 = _GEN_386[26];
          _GEN_122 = _GEN_386[27];
          _GEN_123 = _GEN_386[28];
          _GEN_124 = _GEN_386[29];
          _GEN_125 = _GEN_386[30];
          _GEN_126 = _GEN_386[31];
        end
        else if (inst[31:20] == 12'h321) begin
          _GEN_127 = _GEN_386[0];
          _GEN_128 = _GEN_386[1];
          _GEN_129 = _GEN_386[2];
          _GEN_130 = _GEN_386[3];
          _GEN_131 = _GEN_386[4];
          _GEN_132 = _GEN_386[5];
          _GEN_133 = _GEN_386[6];
          _GEN_134 = _GEN_386[7];
          _GEN_135 = _GEN_386[8];
          _GEN_136 = _GEN_386[9];
          _GEN_137 = _GEN_386[10];
          _GEN_138 = _GEN_386[11];
          _GEN_139 = _GEN_386[12];
          _GEN_140 = _GEN_386[13];
          _GEN_141 = _GEN_386[14];
          _GEN_142 = _GEN_386[15];
          _GEN_143 = _GEN_386[16];
          _GEN_144 = _GEN_386[17];
          _GEN_145 = _GEN_386[18];
          _GEN_146 = _GEN_386[19];
          _GEN_147 = _GEN_386[20];
          _GEN_148 = _GEN_386[21];
          _GEN_149 = _GEN_386[22];
          _GEN_150 = _GEN_386[23];
          _GEN_151 = _GEN_386[24];
          _GEN_152 = _GEN_386[25];
          _GEN_153 = _GEN_386[26];
          _GEN_154 = _GEN_386[27];
          _GEN_155 = _GEN_386[28];
          _GEN_156 = _GEN_386[29];
          _GEN_157 = _GEN_386[30];
          _GEN_158 = _GEN_386[31];
        end
        else if (inst[31:20] == 12'h340) begin
          _GEN_159 = _GEN_386[0];
          _GEN_160 = _GEN_386[1];
          _GEN_161 = _GEN_386[2];
          _GEN_162 = _GEN_386[3];
          _GEN_163 = _GEN_386[4];
          _GEN_164 = _GEN_386[5];
          _GEN_165 = _GEN_386[6];
          _GEN_166 = _GEN_386[7];
          _GEN_167 = _GEN_386[8];
          _GEN_168 = _GEN_386[9];
          _GEN_169 = _GEN_386[10];
          _GEN_170 = _GEN_386[11];
          _GEN_171 = _GEN_386[12];
          _GEN_172 = _GEN_386[13];
          _GEN_173 = _GEN_386[14];
          _GEN_174 = _GEN_386[15];
          _GEN_175 = _GEN_386[16];
          _GEN_176 = _GEN_386[17];
          _GEN_177 = _GEN_386[18];
          _GEN_178 = _GEN_386[19];
          _GEN_179 = _GEN_386[20];
          _GEN_180 = _GEN_386[21];
          _GEN_181 = _GEN_386[22];
          _GEN_182 = _GEN_386[23];
          _GEN_183 = _GEN_386[24];
          _GEN_184 = _GEN_386[25];
          _GEN_185 = _GEN_386[26];
          _GEN_186 = _GEN_386[27];
          _GEN_187 = _GEN_386[28];
          _GEN_188 = _GEN_386[29];
          _GEN_189 = _GEN_386[30];
          _GEN_190 = _GEN_386[31];
        end
        else if (inst[31:20] == 12'h341)
          _GEN_19 = {_GEN_386[31:2], 2'h0};
        else if (inst[31:20] == 12'h342)
          _GEN_20 = _GEN_386 & 32'h8000000F;
        else if (inst[31:20] == 12'h343) begin
          _GEN_27 = _GEN_386[0];
          _GEN_28 = _GEN_386[1];
          _GEN_29 = _GEN_386[2];
          _GEN_30 = _GEN_386[3];
          _GEN_31 = _GEN_386[4];
          _GEN_32 = _GEN_386[5];
          _GEN_33 = _GEN_386[6];
          _GEN_34 = _GEN_386[7];
          _GEN_35 = _GEN_386[8];
          _GEN_36 = _GEN_386[9];
          _GEN_37 = _GEN_386[10];
          _GEN_38 = _GEN_386[11];
          _GEN_39 = _GEN_386[12];
          _GEN_40 = _GEN_386[13];
          _GEN_41 = _GEN_386[14];
          _GEN_42 = _GEN_386[15];
          _GEN_43 = _GEN_386[16];
          _GEN_44 = _GEN_386[17];
          _GEN_45 = _GEN_386[18];
          _GEN_46 = _GEN_386[19];
          _GEN_47 = _GEN_386[20];
          _GEN_48 = _GEN_386[21];
          _GEN_49 = _GEN_386[22];
          _GEN_50 = _GEN_386[23];
          _GEN_51 = _GEN_386[24];
          _GEN_52 = _GEN_386[25];
          _GEN_53 = _GEN_386[26];
          _GEN_54 = _GEN_386[27];
          _GEN_55 = _GEN_386[28];
          _GEN_56 = _GEN_386[29];
          _GEN_57 = _GEN_386[30];
          _GEN_58 = _GEN_386[31];
        end
        else if (inst[31:20] == 12'h780) begin
          _GEN_191 = _GEN_386[0];
          _GEN_192 = _GEN_386[1];
          _GEN_193 = _GEN_386[2];
          _GEN_194 = _GEN_386[3];
          _GEN_195 = _GEN_386[4];
          _GEN_196 = _GEN_386[5];
          _GEN_197 = _GEN_386[6];
          _GEN_198 = _GEN_386[7];
          _GEN_199 = _GEN_386[8];
          _GEN_200 = _GEN_386[9];
          _GEN_201 = _GEN_386[10];
          _GEN_202 = _GEN_386[11];
          _GEN_203 = _GEN_386[12];
          _GEN_204 = _GEN_386[13];
          _GEN_205 = _GEN_386[14];
          _GEN_206 = _GEN_386[15];
          _GEN_207 = _GEN_386[16];
          _GEN_208 = _GEN_386[17];
          _GEN_209 = _GEN_386[18];
          _GEN_210 = _GEN_386[19];
          _GEN_211 = _GEN_386[20];
          _GEN_212 = _GEN_386[21];
          _GEN_213 = _GEN_386[22];
          _GEN_214 = _GEN_386[23];
          _GEN_215 = _GEN_386[24];
          _GEN_216 = _GEN_386[25];
          _GEN_217 = _GEN_386[26];
          _GEN_218 = _GEN_386[27];
          _GEN_219 = _GEN_386[28];
          _GEN_220 = _GEN_386[29];
          _GEN_221 = _GEN_386[30];
          _GEN_222 = _GEN_386[31];
        end
        else if (inst[31:20] == 12'h781) begin
          _GEN_223 = _GEN_386[0];
          _GEN_224 = _GEN_386[1];
          _GEN_225 = _GEN_386[2];
          _GEN_226 = _GEN_386[3];
          _GEN_227 = _GEN_386[4];
          _GEN_228 = _GEN_386[5];
          _GEN_229 = _GEN_386[6];
          _GEN_230 = _GEN_386[7];
          _GEN_231 = _GEN_386[8];
          _GEN_232 = _GEN_386[9];
          _GEN_233 = _GEN_386[10];
          _GEN_234 = _GEN_386[11];
          _GEN_235 = _GEN_386[12];
          _GEN_236 = _GEN_386[13];
          _GEN_237 = _GEN_386[14];
          _GEN_238 = _GEN_386[15];
          _GEN_239 = _GEN_386[16];
          _GEN_240 = _GEN_386[17];
          _GEN_241 = _GEN_386[18];
          _GEN_242 = _GEN_386[19];
          _GEN_243 = _GEN_386[20];
          _GEN_244 = _GEN_386[21];
          _GEN_245 = _GEN_386[22];
          _GEN_246 = _GEN_386[23];
          _GEN_247 = _GEN_386[24];
          _GEN_248 = _GEN_386[25];
          _GEN_249 = _GEN_386[26];
          _GEN_250 = _GEN_386[27];
          _GEN_251 = _GEN_386[28];
          _GEN_252 = _GEN_386[29];
          _GEN_253 = _GEN_386[30];
          _GEN_254 = _GEN_386[31];
        end
        else if (inst[31:20] == 12'h900) begin
          _GEN_255 = _GEN_386[0];
          _GEN_256 = _GEN_386[1];
          _GEN_257 = _GEN_386[2];
          _GEN_258 = _GEN_386[3];
          _GEN_259 = _GEN_386[4];
          _GEN_260 = _GEN_386[5];
          _GEN_261 = _GEN_386[6];
          _GEN_262 = _GEN_386[7];
          _GEN_263 = _GEN_386[8];
          _GEN_264 = _GEN_386[9];
          _GEN_265 = _GEN_386[10];
          _GEN_266 = _GEN_386[11];
          _GEN_267 = _GEN_386[12];
          _GEN_268 = _GEN_386[13];
          _GEN_269 = _GEN_386[14];
          _GEN_270 = _GEN_386[15];
          _GEN_271 = _GEN_386[16];
          _GEN_272 = _GEN_386[17];
          _GEN_273 = _GEN_386[18];
          _GEN_274 = _GEN_386[19];
          _GEN_275 = _GEN_386[20];
          _GEN_276 = _GEN_386[21];
          _GEN_277 = _GEN_386[22];
          _GEN_278 = _GEN_386[23];
          _GEN_279 = _GEN_386[24];
          _GEN_280 = _GEN_386[25];
          _GEN_281 = _GEN_386[26];
          _GEN_282 = _GEN_386[27];
          _GEN_283 = _GEN_386[28];
          _GEN_284 = _GEN_386[29];
          _GEN_285 = _GEN_386[30];
          _GEN_286 = _GEN_386[31];
        end
        else if (inst[31:20] == 12'h901) begin
          _GEN_63 = _GEN_386[0];
          _GEN_64 = _GEN_386[1];
          _GEN_65 = _GEN_386[2];
          _GEN_66 = _GEN_386[3];
          _GEN_67 = _GEN_386[4];
          _GEN_68 = _GEN_386[5];
          _GEN_69 = _GEN_386[6];
          _GEN_70 = _GEN_386[7];
          _GEN_71 = _GEN_386[8];
          _GEN_72 = _GEN_386[9];
          _GEN_73 = _GEN_386[10];
          _GEN_74 = _GEN_386[11];
          _GEN_75 = _GEN_386[12];
          _GEN_76 = _GEN_386[13];
          _GEN_77 = _GEN_386[14];
          _GEN_78 = _GEN_386[15];
          _GEN_79 = _GEN_386[16];
          _GEN_80 = _GEN_386[17];
          _GEN_81 = _GEN_386[18];
          _GEN_82 = _GEN_386[19];
          _GEN_83 = _GEN_386[20];
          _GEN_84 = _GEN_386[21];
          _GEN_85 = _GEN_386[22];
          _GEN_86 = _GEN_386[23];
          _GEN_87 = _GEN_386[24];
          _GEN_88 = _GEN_386[25];
          _GEN_89 = _GEN_386[26];
          _GEN_90 = _GEN_386[27];
          _GEN_91 = _GEN_386[28];
          _GEN_92 = _GEN_386[29];
          _GEN_93 = _GEN_386[30];
          _GEN_94 = _GEN_386[31];
        end
        else if (inst[31:20] == 12'h902) begin
          _GEN_287 = _GEN_386[0];
          _GEN_288 = _GEN_386[1];
          _GEN_289 = _GEN_386[2];
          _GEN_290 = _GEN_386[3];
          _GEN_291 = _GEN_386[4];
          _GEN_292 = _GEN_386[5];
          _GEN_293 = _GEN_386[6];
          _GEN_294 = _GEN_386[7];
          _GEN_295 = _GEN_386[8];
          _GEN_296 = _GEN_386[9];
          _GEN_297 = _GEN_386[10];
          _GEN_298 = _GEN_386[11];
          _GEN_299 = _GEN_386[12];
          _GEN_300 = _GEN_386[13];
          _GEN_301 = _GEN_386[14];
          _GEN_302 = _GEN_386[15];
          _GEN_303 = _GEN_386[16];
          _GEN_304 = _GEN_386[17];
          _GEN_305 = _GEN_386[18];
          _GEN_306 = _GEN_386[19];
          _GEN_307 = _GEN_386[20];
          _GEN_308 = _GEN_386[21];
          _GEN_309 = _GEN_386[22];
          _GEN_310 = _GEN_386[23];
          _GEN_311 = _GEN_386[24];
          _GEN_312 = _GEN_386[25];
          _GEN_313 = _GEN_386[26];
          _GEN_314 = _GEN_386[27];
          _GEN_315 = _GEN_386[28];
          _GEN_316 = _GEN_386[29];
          _GEN_317 = _GEN_386[30];
          _GEN_318 = _GEN_386[31];
        end
        else if (inst[31:20] == 12'h980) begin
          _GEN_319 = _GEN_386[0];
          _GEN_320 = _GEN_386[1];
          _GEN_321 = _GEN_386[2];
          _GEN_322 = _GEN_386[3];
          _GEN_323 = _GEN_386[4];
          _GEN_324 = _GEN_386[5];
          _GEN_325 = _GEN_386[6];
          _GEN_326 = _GEN_386[7];
          _GEN_327 = _GEN_386[8];
          _GEN_328 = _GEN_386[9];
          _GEN_329 = _GEN_386[10];
          _GEN_330 = _GEN_386[11];
          _GEN_331 = _GEN_386[12];
          _GEN_332 = _GEN_386[13];
          _GEN_333 = _GEN_386[14];
          _GEN_334 = _GEN_386[15];
          _GEN_335 = _GEN_386[16];
          _GEN_336 = _GEN_386[17];
          _GEN_337 = _GEN_386[18];
          _GEN_338 = _GEN_386[19];
          _GEN_339 = _GEN_386[20];
          _GEN_340 = _GEN_386[21];
          _GEN_341 = _GEN_386[22];
          _GEN_342 = _GEN_386[23];
          _GEN_343 = _GEN_386[24];
          _GEN_344 = _GEN_386[25];
          _GEN_345 = _GEN_386[26];
          _GEN_346 = _GEN_386[27];
          _GEN_347 = _GEN_386[28];
          _GEN_348 = _GEN_386[29];
          _GEN_349 = _GEN_386[30];
          _GEN_350 = _GEN_386[31];
        end
        else if (inst[31:20] == 12'h981) begin
          _GEN_95 = _GEN_386[0];
          _GEN_96 = _GEN_386[1];
          _GEN_97 = _GEN_386[2];
          _GEN_98 = _GEN_386[3];
          _GEN_99 = _GEN_386[4];
          _GEN_100 = _GEN_386[5];
          _GEN_101 = _GEN_386[6];
          _GEN_102 = _GEN_386[7];
          _GEN_103 = _GEN_386[8];
          _GEN_104 = _GEN_386[9];
          _GEN_105 = _GEN_386[10];
          _GEN_106 = _GEN_386[11];
          _GEN_107 = _GEN_386[12];
          _GEN_108 = _GEN_386[13];
          _GEN_109 = _GEN_386[14];
          _GEN_110 = _GEN_386[15];
          _GEN_111 = _GEN_386[16];
          _GEN_112 = _GEN_386[17];
          _GEN_113 = _GEN_386[18];
          _GEN_114 = _GEN_386[19];
          _GEN_115 = _GEN_386[20];
          _GEN_116 = _GEN_386[21];
          _GEN_117 = _GEN_386[22];
          _GEN_118 = _GEN_386[23];
          _GEN_119 = _GEN_386[24];
          _GEN_120 = _GEN_386[25];
          _GEN_121 = _GEN_386[26];
          _GEN_122 = _GEN_386[27];
          _GEN_123 = _GEN_386[28];
          _GEN_124 = _GEN_386[29];
          _GEN_125 = _GEN_386[30];
          _GEN_126 = _GEN_386[31];
        end
        else if (inst[31:20] == 12'h982) begin
          _GEN_351 = _GEN_386[0];
          _GEN_352 = _GEN_386[1];
          _GEN_353 = _GEN_386[2];
          _GEN_354 = _GEN_386[3];
          _GEN_355 = _GEN_386[4];
          _GEN_356 = _GEN_386[5];
          _GEN_357 = _GEN_386[6];
          _GEN_358 = _GEN_386[7];
          _GEN_359 = _GEN_386[8];
          _GEN_360 = _GEN_386[9];
          _GEN_361 = _GEN_386[10];
          _GEN_362 = _GEN_386[11];
          _GEN_363 = _GEN_386[12];
          _GEN_364 = _GEN_386[13];
          _GEN_365 = _GEN_386[14];
          _GEN_366 = _GEN_386[15];
          _GEN_367 = _GEN_386[16];
          _GEN_368 = _GEN_386[17];
          _GEN_369 = _GEN_386[18];
          _GEN_370 = _GEN_386[19];
          _GEN_371 = _GEN_386[20];
          _GEN_372 = _GEN_386[21];
          _GEN_373 = _GEN_386[22];
          _GEN_374 = _GEN_386[23];
          _GEN_375 = _GEN_386[24];
          _GEN_376 = _GEN_386[25];
          _GEN_377 = _GEN_386[26];
          _GEN_378 = _GEN_386[27];
          _GEN_379 = _GEN_386[28];
          _GEN_380 = _GEN_386[29];
          _GEN_381 = _GEN_386[30];
          _GEN_382 = _GEN_386[31];
        end
      end
    end
  end // always_comb
  always_ff @(posedge CLK) begin
    if (RESET) begin
      Register_inst6 <= 2'h3;
      Register_inst16 <= 32'h0;
      Register_inst17 <= 32'h0;
      Register_inst8 <= 1'h0;
      Register_inst7 <= 2'h3;
      Register_inst9 <= 1'h0;
      Register_inst18 <= 32'h0;
      Register_inst10 <= 1'h0;
      Register_inst12 <= 1'h0;
      Register_inst11 <= 1'h0;
      Register_inst13 <= 1'h0;
      Register_inst0 <= 32'h0;
      Register_inst1 <= 32'h0;
      Register_inst14 <= 32'h0;
      Register_inst15 <= 32'h0;
      Register_inst19 <= 32'h0;
      Register_inst20 <= 32'h0;
      Register_inst4 <= 32'h0;
      Register_inst3 <= 32'h0;
      Register_inst5 <= 32'h0;
      Register_inst2 <= 32'h0;
    end
    else begin
      Register_inst6 <= {_GEN_22, _GEN_21};
      Register_inst16 <= _GEN_19;
      Register_inst17 <= _GEN_20;
      Register_inst8 <= _GEN_23;
      Register_inst7 <= {_GEN_25, _GEN_24};
      Register_inst9 <= _GEN_26;
      Register_inst18 <=
        {_GEN_58,
         _GEN_57,
         _GEN_56,
         _GEN_55,
         _GEN_54,
         _GEN_53,
         _GEN_52,
         _GEN_51,
         _GEN_50,
         _GEN_49,
         _GEN_48,
         _GEN_47,
         _GEN_46,
         _GEN_45,
         _GEN_44,
         _GEN_43,
         _GEN_42,
         _GEN_41,
         _GEN_40,
         _GEN_39,
         _GEN_38,
         _GEN_37,
         _GEN_36,
         _GEN_35,
         _GEN_34,
         _GEN_33,
         _GEN_32,
         _GEN_31,
         _GEN_30,
         _GEN_29,
         _GEN_28,
         _GEN_27};
      Register_inst10 <= _GEN_59;
      Register_inst12 <= _GEN_60;
      Register_inst11 <= _GEN_61;
      Register_inst13 <= _GEN_62;
      Register_inst0 <=
        {_GEN_94,
         _GEN_93,
         _GEN_92,
         _GEN_91,
         _GEN_90,
         _GEN_89,
         _GEN_88,
         _GEN_87,
         _GEN_86,
         _GEN_85,
         _GEN_84,
         _GEN_83,
         _GEN_82,
         _GEN_81,
         _GEN_80,
         _GEN_79,
         _GEN_78,
         _GEN_77,
         _GEN_76,
         _GEN_75,
         _GEN_74,
         _GEN_73,
         _GEN_72,
         _GEN_71,
         _GEN_70,
         _GEN_69,
         _GEN_68,
         _GEN_67,
         _GEN_66,
         _GEN_65,
         _GEN_64,
         _GEN_63};
      Register_inst1 <=
        {_GEN_126,
         _GEN_125,
         _GEN_124,
         _GEN_123,
         _GEN_122,
         _GEN_121,
         _GEN_120,
         _GEN_119,
         _GEN_118,
         _GEN_117,
         _GEN_116,
         _GEN_115,
         _GEN_114,
         _GEN_113,
         _GEN_112,
         _GEN_111,
         _GEN_110,
         _GEN_109,
         _GEN_108,
         _GEN_107,
         _GEN_106,
         _GEN_105,
         _GEN_104,
         _GEN_103,
         _GEN_102,
         _GEN_101,
         _GEN_100,
         _GEN_99,
         _GEN_98,
         _GEN_97,
         _GEN_96,
         _GEN_95};
      Register_inst14 <=
        {_GEN_158,
         _GEN_157,
         _GEN_156,
         _GEN_155,
         _GEN_154,
         _GEN_153,
         _GEN_152,
         _GEN_151,
         _GEN_150,
         _GEN_149,
         _GEN_148,
         _GEN_147,
         _GEN_146,
         _GEN_145,
         _GEN_144,
         _GEN_143,
         _GEN_142,
         _GEN_141,
         _GEN_140,
         _GEN_139,
         _GEN_138,
         _GEN_137,
         _GEN_136,
         _GEN_135,
         _GEN_134,
         _GEN_133,
         _GEN_132,
         _GEN_131,
         _GEN_130,
         _GEN_129,
         _GEN_128,
         _GEN_127};
      Register_inst15 <=
        {_GEN_190,
         _GEN_189,
         _GEN_188,
         _GEN_187,
         _GEN_186,
         _GEN_185,
         _GEN_184,
         _GEN_183,
         _GEN_182,
         _GEN_181,
         _GEN_180,
         _GEN_179,
         _GEN_178,
         _GEN_177,
         _GEN_176,
         _GEN_175,
         _GEN_174,
         _GEN_173,
         _GEN_172,
         _GEN_171,
         _GEN_170,
         _GEN_169,
         _GEN_168,
         _GEN_167,
         _GEN_166,
         _GEN_165,
         _GEN_164,
         _GEN_163,
         _GEN_162,
         _GEN_161,
         _GEN_160,
         _GEN_159};
      Register_inst19 <=
        {_GEN_222,
         _GEN_221,
         _GEN_220,
         _GEN_219,
         _GEN_218,
         _GEN_217,
         _GEN_216,
         _GEN_215,
         _GEN_214,
         _GEN_213,
         _GEN_212,
         _GEN_211,
         _GEN_210,
         _GEN_209,
         _GEN_208,
         _GEN_207,
         _GEN_206,
         _GEN_205,
         _GEN_204,
         _GEN_203,
         _GEN_202,
         _GEN_201,
         _GEN_200,
         _GEN_199,
         _GEN_198,
         _GEN_197,
         _GEN_196,
         _GEN_195,
         _GEN_194,
         _GEN_193,
         _GEN_192,
         _GEN_191};
      Register_inst20 <=
        {_GEN_254,
         _GEN_253,
         _GEN_252,
         _GEN_251,
         _GEN_250,
         _GEN_249,
         _GEN_248,
         _GEN_247,
         _GEN_246,
         _GEN_245,
         _GEN_244,
         _GEN_243,
         _GEN_242,
         _GEN_241,
         _GEN_240,
         _GEN_239,
         _GEN_238,
         _GEN_237,
         _GEN_236,
         _GEN_235,
         _GEN_234,
         _GEN_233,
         _GEN_232,
         _GEN_231,
         _GEN_230,
         _GEN_229,
         _GEN_228,
         _GEN_227,
         _GEN_226,
         _GEN_225,
         _GEN_224,
         _GEN_223};
      Register_inst4 <=
        {_GEN_318,
         _GEN_317,
         _GEN_316,
         _GEN_315,
         _GEN_314,
         _GEN_313,
         _GEN_312,
         _GEN_311,
         _GEN_310,
         _GEN_309,
         _GEN_308,
         _GEN_307,
         _GEN_306,
         _GEN_305,
         _GEN_304,
         _GEN_303,
         _GEN_302,
         _GEN_301,
         _GEN_300,
         _GEN_299,
         _GEN_298,
         _GEN_297,
         _GEN_296,
         _GEN_295,
         _GEN_294,
         _GEN_293,
         _GEN_292,
         _GEN_291,
         _GEN_290,
         _GEN_289,
         _GEN_288,
         _GEN_287};
      Register_inst3 <=
        {_GEN_350,
         _GEN_349,
         _GEN_348,
         _GEN_347,
         _GEN_346,
         _GEN_345,
         _GEN_344,
         _GEN_343,
         _GEN_342,
         _GEN_341,
         _GEN_340,
         _GEN_339,
         _GEN_338,
         _GEN_337,
         _GEN_336,
         _GEN_335,
         _GEN_334,
         _GEN_333,
         _GEN_332,
         _GEN_331,
         _GEN_330,
         _GEN_329,
         _GEN_328,
         _GEN_327,
         _GEN_326,
         _GEN_325,
         _GEN_324,
         _GEN_323,
         _GEN_322,
         _GEN_321,
         _GEN_320,
         _GEN_319};
      Register_inst5 <=
        {_GEN_382,
         _GEN_381,
         _GEN_380,
         _GEN_379,
         _GEN_378,
         _GEN_377,
         _GEN_376,
         _GEN_375,
         _GEN_374,
         _GEN_373,
         _GEN_372,
         _GEN_371,
         _GEN_370,
         _GEN_369,
         _GEN_368,
         _GEN_367,
         _GEN_366,
         _GEN_365,
         _GEN_364,
         _GEN_363,
         _GEN_362,
         _GEN_361,
         _GEN_360,
         _GEN_359,
         _GEN_358,
         _GEN_357,
         _GEN_356,
         _GEN_355,
         _GEN_354,
         _GEN_353,
         _GEN_352,
         _GEN_351};
      Register_inst2 <=
        {_GEN_286,
         _GEN_285,
         _GEN_284,
         _GEN_283,
         _GEN_282,
         _GEN_281,
         _GEN_280,
         _GEN_279,
         _GEN_278,
         _GEN_277,
         _GEN_276,
         _GEN_275,
         _GEN_274,
         _GEN_273,
         _GEN_272,
         _GEN_271,
         _GEN_270,
         _GEN_269,
         _GEN_268,
         _GEN_267,
         _GEN_266,
         _GEN_265,
         _GEN_264,
         _GEN_263,
         _GEN_262,
         _GEN_261,
         _GEN_260,
         _GEN_259,
         _GEN_258,
         _GEN_257,
         _GEN_256,
         _GEN_255};
    end
  end // always_ff @(posedge)
  initial begin
    Register_inst6 = 2'h3;
    Register_inst16 = 32'h0;
    Register_inst17 = 32'h0;
    Register_inst8 = 1'h0;
    Register_inst7 = 2'h3;
    Register_inst9 = 1'h0;
    Register_inst18 = 32'h0;
    Register_inst10 = 1'h0;
    Register_inst12 = 1'h0;
    Register_inst11 = 1'h0;
    Register_inst13 = 1'h0;
    Register_inst0 = 32'h0;
    Register_inst1 = 32'h0;
    Register_inst14 = 32'h0;
    Register_inst15 = 32'h0;
    Register_inst19 = 32'h0;
    Register_inst20 = 32'h0;
    Register_inst4 = 32'h0;
    Register_inst3 = 32'h0;
    Register_inst5 = 32'h0;
    Register_inst2 = 32'h0;
  end // initial
  wire [1:0][31:0] _GEN_389 = {{Register_inst2}, {32'h0}};
  wire [1:0][31:0] _GEN_390 = {{Register_inst0}, {_GEN_389[inst[31:20] == 12'hC00]}};
  wire [1:0][31:0] _GEN_391 = {{Register_inst4}, {_GEN_390[inst[31:20] == 12'hC01]}};
  wire [1:0][31:0] _GEN_392 = {{Register_inst3}, {_GEN_391[inst[31:20] == 12'hC02]}};
  wire [1:0][31:0] _GEN_393 = {{Register_inst1}, {_GEN_392[inst[31:20] == 12'hC80]}};
  wire [1:0][31:0] _GEN_394 = {{Register_inst5}, {_GEN_393[inst[31:20] == 12'hC81]}};
  wire [1:0][31:0] _GEN_395 = {{Register_inst2}, {_GEN_394[inst[31:20] == 12'hC82]}};
  wire [1:0][31:0] _GEN_396 = {{Register_inst0}, {_GEN_395[inst[31:20] == 12'h900]}};
  wire [1:0][31:0] _GEN_397 = {{Register_inst4}, {_GEN_396[inst[31:20] == 12'h901]}};
  wire [1:0][31:0] _GEN_398 = {{Register_inst3}, {_GEN_397[inst[31:20] == 12'h902]}};
  wire [1:0][31:0] _GEN_399 = {{Register_inst1}, {_GEN_398[inst[31:20] == 12'h980]}};
  wire [1:0][31:0] _GEN_400 = {{Register_inst5}, {_GEN_399[inst[31:20] == 12'h981]}};
  wire [1:0][31:0] _GEN_401 = {{32'h100100}, {_GEN_400[inst[31:20] == 12'h982]}};
  wire [1:0][31:0] _GEN_402 = {{32'h0}, {_GEN_401[inst[31:20] == 12'hF00]}};
  wire [1:0][31:0] _GEN_403 = {{32'h0}, {_GEN_402[inst[31:20] == 12'hF01]}};
  wire [1:0][31:0] _GEN_404 = {{32'h100}, {_GEN_403[inst[31:20] == 12'hF10]}};
  wire [1:0][31:0] _GEN_405 = {{32'h0}, {_GEN_404[inst[31:20] == 12'h301]}};
  wire [1:0][31:0] _GEN_406 =
    {{{24'h0, Register_inst11, 3'h0, Register_inst13, 3'h0}},
     {_GEN_405[inst[31:20] == 12'h302]}};
  wire [1:0][31:0] _GEN_407 = {{Register_inst14}, {_GEN_406[inst[31:20] == 12'h304]}};
  wire [1:0][31:0] _GEN_408 = {{Register_inst0}, {_GEN_407[inst[31:20] == 12'h321]}};
  wire [1:0][31:0] _GEN_409 = {{Register_inst1}, {_GEN_408[inst[31:20] == 12'h701]}};
  wire [1:0][31:0] _GEN_410 = {{Register_inst15}, {_GEN_409[inst[31:20] == 12'h741]}};
  wire [1:0][31:0] _GEN_411 = {{Register_inst16}, {_GEN_410[inst[31:20] == 12'h340]}};
  wire [1:0][31:0] _GEN_412 = {{Register_inst17}, {_GEN_411[inst[31:20] == 12'h341]}};
  wire [1:0][31:0] _GEN_413 = {{Register_inst18}, {_GEN_412[inst[31:20] == 12'h342]}};
  wire [1:0][31:0] _GEN_414 =
    {{{24'h0, Register_inst10, 3'h0, Register_inst12, 3'h0}},
     {_GEN_413[inst[31:20] == 12'h343]}};
  wire [1:0][31:0] _GEN_415 = {{Register_inst19}, {_GEN_414[inst[31:20] == 12'h344]}};
  wire [1:0][31:0] _GEN_416 = {{Register_inst20}, {_GEN_415[inst[31:20] == 12'h780]}};
  wire [1:0][31:0] _GEN_417 =
    {{{26'h0, Register_inst7, Register_inst9, Register_inst6, Register_inst8}},
     {_GEN_416[inst[31:20] == 12'h781]}};
  assign _GEN = _GEN_417[inst[31:20] == 12'h300];
  assign O = _GEN;
  assign expt = _GEN_13;
  assign evec = {24'h0, Register_inst6, 6'h0} + 32'h100;
  assign epc = Register_inst16;
  assign host_tohost = Register_inst19;
endmodule

module RegFile(
  input  [4:0]  raddr1,
                raddr2,
  input         wen,
  input  [4:0]  waddr,
  input  [31:0] wdata,
  input         CLK,
                RESET,
  output [31:0] rdata1,
                rdata2
);

  reg  [31:0][31:0] MultiportMemory_inst0;
  always_ff @(posedge CLK) begin
    if (wen & (|waddr))
      MultiportMemory_inst0[waddr] <= wdata;
  end // always_ff @(posedge)
  wire [1:0][31:0]  _GEN = {{MultiportMemory_inst0[raddr1]}, {32'h0}};
  wire [1:0][31:0]  _GEN_0 = {{MultiportMemory_inst0[raddr2]}, {32'h0}};
  assign rdata1 = _GEN[|raddr1];
  assign rdata2 = _GEN_0[|raddr2];
endmodule

module ALUArea(
  input  [31:0] A,
                B,
  input  [3:0]  op,
  output [31:0] O,
                sum_
);

  wire [1:0][31:0] _GEN = {{32'h0 - B}, {B}};
  wire [31:0]      _GEN_0 = A + _GEN[op[0]];
  reg              _GEN_1;
  reg              _GEN_2;
  reg              _GEN_3;
  reg              _GEN_4;
  reg              _GEN_5;
  reg              _GEN_6;
  reg              _GEN_7;
  reg              _GEN_8;
  reg              _GEN_9;
  reg              _GEN_10;
  reg              _GEN_11;
  reg              _GEN_12;
  reg              _GEN_13;
  reg              _GEN_14;
  reg              _GEN_15;
  reg              _GEN_16;
  reg              _GEN_17;
  reg              _GEN_18;
  reg              _GEN_19;
  reg              _GEN_20;
  reg              _GEN_21;
  reg              _GEN_22;
  reg              _GEN_23;
  reg              _GEN_24;
  reg              _GEN_25;
  reg              _GEN_26;
  reg              _GEN_27;
  reg              _GEN_28;
  reg              _GEN_29;
  reg              _GEN_30;
  reg              _GEN_31;
  reg              _GEN_32;
  wire [31:0]      _GEN_33 = A & B;
  wire [31:0]      _GEN_34 = A | B;
  wire [31:0]      _GEN_35 = A ^ B;
  wire [1:0]       _GEN_36 = {{B[31]}, {A[31]}};
  wire [1:0][31:0] _GEN_37 =
    {{A},
     {{A[0],
       A[1],
       A[2],
       A[3],
       A[4],
       A[5],
       A[6],
       A[7],
       A[8],
       A[9],
       A[10],
       A[11],
       A[12],
       A[13],
       A[14],
       A[15],
       A[16],
       A[17],
       A[18],
       A[19],
       A[20],
       A[21],
       A[22],
       A[23],
       A[24],
       A[25],
       A[26],
       A[27],
       A[28],
       A[29],
       A[30],
       A[31]}}};
  wire [31:0]      _GEN_38 = _GEN_37[op[3]];
  wire [32:0]      _GEN_39 = $signed($signed({op[0] & _GEN_38[31], _GEN_38}) >>> B);
  wire [1:0]       _GEN_40 = {{_GEN_0[31]}, {_GEN_36[op[1]]}};
  always_comb begin
    if (op == 4'h0 | op == 4'h1) begin
      _GEN_1 = _GEN_0[0];
      _GEN_2 = _GEN_0[1];
      _GEN_3 = _GEN_0[2];
      _GEN_4 = _GEN_0[3];
      _GEN_5 = _GEN_0[4];
      _GEN_6 = _GEN_0[5];
      _GEN_7 = _GEN_0[6];
      _GEN_8 = _GEN_0[7];
      _GEN_9 = _GEN_0[8];
      _GEN_10 = _GEN_0[9];
      _GEN_11 = _GEN_0[10];
      _GEN_12 = _GEN_0[11];
      _GEN_13 = _GEN_0[12];
      _GEN_14 = _GEN_0[13];
      _GEN_15 = _GEN_0[14];
      _GEN_16 = _GEN_0[15];
      _GEN_17 = _GEN_0[16];
      _GEN_18 = _GEN_0[17];
      _GEN_19 = _GEN_0[18];
      _GEN_20 = _GEN_0[19];
      _GEN_21 = _GEN_0[20];
      _GEN_22 = _GEN_0[21];
      _GEN_23 = _GEN_0[22];
      _GEN_24 = _GEN_0[23];
      _GEN_25 = _GEN_0[24];
      _GEN_26 = _GEN_0[25];
      _GEN_27 = _GEN_0[26];
      _GEN_28 = _GEN_0[27];
      _GEN_29 = _GEN_0[28];
      _GEN_30 = _GEN_0[29];
      _GEN_31 = _GEN_0[30];
      _GEN_32 = _GEN_0[31];
    end
    else if (op == 4'h5 | op == 4'h7) begin
      _GEN_1 = _GEN_40[A[31] ^ ~(B[31])];
      _GEN_2 = 1'h0;
      _GEN_3 = 1'h0;
      _GEN_4 = 1'h0;
      _GEN_5 = 1'h0;
      _GEN_6 = 1'h0;
      _GEN_7 = 1'h0;
      _GEN_8 = 1'h0;
      _GEN_9 = 1'h0;
      _GEN_10 = 1'h0;
      _GEN_11 = 1'h0;
      _GEN_12 = 1'h0;
      _GEN_13 = 1'h0;
      _GEN_14 = 1'h0;
      _GEN_15 = 1'h0;
      _GEN_16 = 1'h0;
      _GEN_17 = 1'h0;
      _GEN_18 = 1'h0;
      _GEN_19 = 1'h0;
      _GEN_20 = 1'h0;
      _GEN_21 = 1'h0;
      _GEN_22 = 1'h0;
      _GEN_23 = 1'h0;
      _GEN_24 = 1'h0;
      _GEN_25 = 1'h0;
      _GEN_26 = 1'h0;
      _GEN_27 = 1'h0;
      _GEN_28 = 1'h0;
      _GEN_29 = 1'h0;
      _GEN_30 = 1'h0;
      _GEN_31 = 1'h0;
      _GEN_32 = 1'h0;
    end
    else if (op == 4'h9 | op == 4'h8) begin
      _GEN_1 = _GEN_39[0];
      _GEN_2 = _GEN_39[1];
      _GEN_3 = _GEN_39[2];
      _GEN_4 = _GEN_39[3];
      _GEN_5 = _GEN_39[4];
      _GEN_6 = _GEN_39[5];
      _GEN_7 = _GEN_39[6];
      _GEN_8 = _GEN_39[7];
      _GEN_9 = _GEN_39[8];
      _GEN_10 = _GEN_39[9];
      _GEN_11 = _GEN_39[10];
      _GEN_12 = _GEN_39[11];
      _GEN_13 = _GEN_39[12];
      _GEN_14 = _GEN_39[13];
      _GEN_15 = _GEN_39[14];
      _GEN_16 = _GEN_39[15];
      _GEN_17 = _GEN_39[16];
      _GEN_18 = _GEN_39[17];
      _GEN_19 = _GEN_39[18];
      _GEN_20 = _GEN_39[19];
      _GEN_21 = _GEN_39[20];
      _GEN_22 = _GEN_39[21];
      _GEN_23 = _GEN_39[22];
      _GEN_24 = _GEN_39[23];
      _GEN_25 = _GEN_39[24];
      _GEN_26 = _GEN_39[25];
      _GEN_27 = _GEN_39[26];
      _GEN_28 = _GEN_39[27];
      _GEN_29 = _GEN_39[28];
      _GEN_30 = _GEN_39[29];
      _GEN_31 = _GEN_39[30];
      _GEN_32 = _GEN_39[31];
    end
    else if (op == 4'h6) begin
      _GEN_1 = _GEN_39[31];
      _GEN_2 = _GEN_39[30];
      _GEN_3 = _GEN_39[29];
      _GEN_4 = _GEN_39[28];
      _GEN_5 = _GEN_39[27];
      _GEN_6 = _GEN_39[26];
      _GEN_7 = _GEN_39[25];
      _GEN_8 = _GEN_39[24];
      _GEN_9 = _GEN_39[23];
      _GEN_10 = _GEN_39[22];
      _GEN_11 = _GEN_39[21];
      _GEN_12 = _GEN_39[20];
      _GEN_13 = _GEN_39[19];
      _GEN_14 = _GEN_39[18];
      _GEN_15 = _GEN_39[17];
      _GEN_16 = _GEN_39[16];
      _GEN_17 = _GEN_39[15];
      _GEN_18 = _GEN_39[14];
      _GEN_19 = _GEN_39[13];
      _GEN_20 = _GEN_39[12];
      _GEN_21 = _GEN_39[11];
      _GEN_22 = _GEN_39[10];
      _GEN_23 = _GEN_39[9];
      _GEN_24 = _GEN_39[8];
      _GEN_25 = _GEN_39[7];
      _GEN_26 = _GEN_39[6];
      _GEN_27 = _GEN_39[5];
      _GEN_28 = _GEN_39[4];
      _GEN_29 = _GEN_39[3];
      _GEN_30 = _GEN_39[2];
      _GEN_31 = _GEN_39[1];
      _GEN_32 = _GEN_39[0];
    end
    else if (op == 4'h2) begin
      _GEN_1 = _GEN_33[0];
      _GEN_2 = _GEN_33[1];
      _GEN_3 = _GEN_33[2];
      _GEN_4 = _GEN_33[3];
      _GEN_5 = _GEN_33[4];
      _GEN_6 = _GEN_33[5];
      _GEN_7 = _GEN_33[6];
      _GEN_8 = _GEN_33[7];
      _GEN_9 = _GEN_33[8];
      _GEN_10 = _GEN_33[9];
      _GEN_11 = _GEN_33[10];
      _GEN_12 = _GEN_33[11];
      _GEN_13 = _GEN_33[12];
      _GEN_14 = _GEN_33[13];
      _GEN_15 = _GEN_33[14];
      _GEN_16 = _GEN_33[15];
      _GEN_17 = _GEN_33[16];
      _GEN_18 = _GEN_33[17];
      _GEN_19 = _GEN_33[18];
      _GEN_20 = _GEN_33[19];
      _GEN_21 = _GEN_33[20];
      _GEN_22 = _GEN_33[21];
      _GEN_23 = _GEN_33[22];
      _GEN_24 = _GEN_33[23];
      _GEN_25 = _GEN_33[24];
      _GEN_26 = _GEN_33[25];
      _GEN_27 = _GEN_33[26];
      _GEN_28 = _GEN_33[27];
      _GEN_29 = _GEN_33[28];
      _GEN_30 = _GEN_33[29];
      _GEN_31 = _GEN_33[30];
      _GEN_32 = _GEN_33[31];
    end
    else if (op == 4'h3) begin
      _GEN_1 = _GEN_34[0];
      _GEN_2 = _GEN_34[1];
      _GEN_3 = _GEN_34[2];
      _GEN_4 = _GEN_34[3];
      _GEN_5 = _GEN_34[4];
      _GEN_6 = _GEN_34[5];
      _GEN_7 = _GEN_34[6];
      _GEN_8 = _GEN_34[7];
      _GEN_9 = _GEN_34[8];
      _GEN_10 = _GEN_34[9];
      _GEN_11 = _GEN_34[10];
      _GEN_12 = _GEN_34[11];
      _GEN_13 = _GEN_34[12];
      _GEN_14 = _GEN_34[13];
      _GEN_15 = _GEN_34[14];
      _GEN_16 = _GEN_34[15];
      _GEN_17 = _GEN_34[16];
      _GEN_18 = _GEN_34[17];
      _GEN_19 = _GEN_34[18];
      _GEN_20 = _GEN_34[19];
      _GEN_21 = _GEN_34[20];
      _GEN_22 = _GEN_34[21];
      _GEN_23 = _GEN_34[22];
      _GEN_24 = _GEN_34[23];
      _GEN_25 = _GEN_34[24];
      _GEN_26 = _GEN_34[25];
      _GEN_27 = _GEN_34[26];
      _GEN_28 = _GEN_34[27];
      _GEN_29 = _GEN_34[28];
      _GEN_30 = _GEN_34[29];
      _GEN_31 = _GEN_34[30];
      _GEN_32 = _GEN_34[31];
    end
    else if (op == 4'h4) begin
      _GEN_1 = _GEN_35[0];
      _GEN_2 = _GEN_35[1];
      _GEN_3 = _GEN_35[2];
      _GEN_4 = _GEN_35[3];
      _GEN_5 = _GEN_35[4];
      _GEN_6 = _GEN_35[5];
      _GEN_7 = _GEN_35[6];
      _GEN_8 = _GEN_35[7];
      _GEN_9 = _GEN_35[8];
      _GEN_10 = _GEN_35[9];
      _GEN_11 = _GEN_35[10];
      _GEN_12 = _GEN_35[11];
      _GEN_13 = _GEN_35[12];
      _GEN_14 = _GEN_35[13];
      _GEN_15 = _GEN_35[14];
      _GEN_16 = _GEN_35[15];
      _GEN_17 = _GEN_35[16];
      _GEN_18 = _GEN_35[17];
      _GEN_19 = _GEN_35[18];
      _GEN_20 = _GEN_35[19];
      _GEN_21 = _GEN_35[20];
      _GEN_22 = _GEN_35[21];
      _GEN_23 = _GEN_35[22];
      _GEN_24 = _GEN_35[23];
      _GEN_25 = _GEN_35[24];
      _GEN_26 = _GEN_35[25];
      _GEN_27 = _GEN_35[26];
      _GEN_28 = _GEN_35[27];
      _GEN_29 = _GEN_35[28];
      _GEN_30 = _GEN_35[29];
      _GEN_31 = _GEN_35[30];
      _GEN_32 = _GEN_35[31];
    end
    else if (op == 4'hA) begin
      _GEN_1 = A[0];
      _GEN_2 = A[1];
      _GEN_3 = A[2];
      _GEN_4 = A[3];
      _GEN_5 = A[4];
      _GEN_6 = A[5];
      _GEN_7 = A[6];
      _GEN_8 = A[7];
      _GEN_9 = A[8];
      _GEN_10 = A[9];
      _GEN_11 = A[10];
      _GEN_12 = A[11];
      _GEN_13 = A[12];
      _GEN_14 = A[13];
      _GEN_15 = A[14];
      _GEN_16 = A[15];
      _GEN_17 = A[16];
      _GEN_18 = A[17];
      _GEN_19 = A[18];
      _GEN_20 = A[19];
      _GEN_21 = A[20];
      _GEN_22 = A[21];
      _GEN_23 = A[22];
      _GEN_24 = A[23];
      _GEN_25 = A[24];
      _GEN_26 = A[25];
      _GEN_27 = A[26];
      _GEN_28 = A[27];
      _GEN_29 = A[28];
      _GEN_30 = A[29];
      _GEN_31 = A[30];
      _GEN_32 = A[31];
    end
    else begin
      _GEN_1 = B[0];
      _GEN_2 = B[1];
      _GEN_3 = B[2];
      _GEN_4 = B[3];
      _GEN_5 = B[4];
      _GEN_6 = B[5];
      _GEN_7 = B[6];
      _GEN_8 = B[7];
      _GEN_9 = B[8];
      _GEN_10 = B[9];
      _GEN_11 = B[10];
      _GEN_12 = B[11];
      _GEN_13 = B[12];
      _GEN_14 = B[13];
      _GEN_15 = B[14];
      _GEN_16 = B[15];
      _GEN_17 = B[16];
      _GEN_18 = B[17];
      _GEN_19 = B[18];
      _GEN_20 = B[19];
      _GEN_21 = B[20];
      _GEN_22 = B[21];
      _GEN_23 = B[22];
      _GEN_24 = B[23];
      _GEN_25 = B[24];
      _GEN_26 = B[25];
      _GEN_27 = B[26];
      _GEN_28 = B[27];
      _GEN_29 = B[28];
      _GEN_30 = B[29];
      _GEN_31 = B[30];
      _GEN_32 = B[31];
    end
  end // always_comb
  assign O =
    {_GEN_32,
     _GEN_31,
     _GEN_30,
     _GEN_29,
     _GEN_28,
     _GEN_27,
     _GEN_26,
     _GEN_25,
     _GEN_24,
     _GEN_23,
     _GEN_22,
     _GEN_21,
     _GEN_20,
     _GEN_19,
     _GEN_18,
     _GEN_17,
     _GEN_16,
     _GEN_15,
     _GEN_14,
     _GEN_13,
     _GEN_12,
     _GEN_11,
     _GEN_10,
     _GEN_9,
     _GEN_8,
     _GEN_7,
     _GEN_6,
     _GEN_5,
     _GEN_4,
     _GEN_3,
     _GEN_2,
     _GEN_1};
  assign sum_ = _GEN_0;
endmodule

module ImmGenWire(
  input  [31:0] inst,
  input  [2:0]  sel,
  output [31:0] O
);

  wire [1:0][31:0] _GEN =
    {{{{21{inst[31]}}, inst[30:20]}}, {{{21{inst[31]}}, inst[30:20]} & 32'hFFFFFFFE}};
  wire [1:0][31:0] _GEN_0 =
    {{{{21{inst[31]}}, inst[30:25], inst[11:7]}}, {_GEN[sel == 3'h1]}};
  wire [1:0][31:0] _GEN_1 =
    {{{{20{inst[31]}}, inst[7], inst[30:25], inst[11:8], 1'h0}}, {_GEN_0[sel == 3'h2]}};
  wire [1:0][31:0] _GEN_2 = {{{inst[31:12], 12'h0}}, {_GEN_1[sel == 3'h5]}};
  wire [1:0][31:0] _GEN_3 =
    {{{{12{inst[31]}}, inst[19:12], inst[20], inst[30:21], 1'h0}}, {_GEN_2[sel == 3'h3]}};
  wire [1:0][31:0] _GEN_4 = {{{27'h0, inst[19:15]}}, {_GEN_3[sel == 3'h4]}};
  assign O = _GEN_4[sel == 3'h6];
endmodule

module BrCondArea(
  input  [31:0] rs1,
                rs2,
  input  [2:0]  br_type,
  output        taken
);

  wire [31:0] _GEN = rs1 - rs2;
  wire        _GEN_0 = rs1[31] ^ ~(rs2[31]);
  wire [1:0]  _GEN_1 = {{_GEN[31]}, {rs1[31]}};
  wire [1:0]  _GEN_2 = {{_GEN[31]}, {rs2[31]}};
  assign taken =
    br_type == 3'h3 & ~(|_GEN) | br_type == 3'h6 & (|_GEN) | br_type == 3'h2
    & _GEN_1[_GEN_0] | br_type == 3'h5 & ~_GEN_1[_GEN_0] | br_type == 3'h1
    & _GEN_2[_GEN_0] | br_type == 3'h4 & ~_GEN_2[_GEN_0];
endmodule

module Datapath(
  input  struct packed {logic valid; logic [31:0] data; }                                                             host_fromhost,
  input  struct packed {logic valid; struct packed {logic [31:0] data; } data; }                                      icache_resp,
                                                                                                                      dcache_resp,
  input  [1:0]                                                                                                        ctrl_pc_sel,
  input                                                                                                               ctrl_inst_kill,
                                                                                                                      ctrl_A_sel,
                                                                                                                      ctrl_B_sel,
  input  [2:0]                                                                                                        ctrl_imm_sel,
  input  [3:0]                                                                                                        ctrl_alu_op,
  input  [2:0]                                                                                                        ctrl_br_type,
  input  [1:0]                                                                                                        ctrl_st_type,
  input  [2:0]                                                                                                        ctrl_ld_type,
  input  [1:0]                                                                                                        ctrl_wb_sel,
  input                                                                                                               ctrl_wb_en,
  input  [2:0]                                                                                                        ctrl_csr_cmd,
  input                                                                                                               ctrl_illegal,
                                                                                                                      CLK,
                                                                                                                      RESET,
  output [31:0]                                                                                                       host_tohost,
  output                                                                                                              icache_abort,
  output struct packed {logic valid; struct packed {logic [31:0] addr; logic [31:0] data; logic [3:0] mask; } data; } icache_req,
  output                                                                                                              dcache_abort,
  output struct packed {logic valid; struct packed {logic [31:0] addr; logic [31:0] data; logic [3:0] mask; } data; } dcache_req,
  output [31:0]                                                                                                       ctrl_inst
);

  reg  [2:0]       Register_inst10;
  reg              _GEN;
  reg              _GEN_0;
  reg              _GEN_1;
  reg              _GEN_2;
  reg              _GEN_3;
  reg              _GEN_4;
  reg              _GEN_5;
  reg              _GEN_6;
  reg              _GEN_7;
  reg              _GEN_8;
  reg              _GEN_9;
  reg              _GEN_10;
  reg              _GEN_11;
  reg              _GEN_12;
  reg              _GEN_13;
  reg              _GEN_14;
  reg              _GEN_15;
  reg              _GEN_16;
  reg              _GEN_17;
  reg              _GEN_18;
  reg              _GEN_19;
  reg              _GEN_20;
  reg              _GEN_21;
  reg              _GEN_22;
  reg              _GEN_23;
  reg              _GEN_24;
  reg              _GEN_25;
  reg              _GEN_26;
  reg              _GEN_27;
  reg              _GEN_28;
  reg              _GEN_29;
  reg              _GEN_30;
  reg  [31:0]      Register_inst1;
  reg  [31:0]      Register_inst14;
  reg  [31:0]      Register_inst0;
  wire [31:0]      _CSRGen_inst0_O;
  wire             _CSRGen_inst0_expt;
  wire [31:0]      _CSRGen_inst0_evec;
  wire [31:0]      _CSRGen_inst0_epc;
  wire [31:0]      _ALUArea_inst0_O;
  wire [31:0]      _ALUArea_inst0_sum_;
  wire [31:0]      _ImmGenWire_inst0_O;
  wire [31:0]      _RegFile_inst0_rdata1;
  wire [31:0]      _RegFile_inst0_rdata2;
  wire             _BrCondArea_inst0_taken;
  wire [1:0][3:0]  _GEN_31 = {4'hF, 4'h0};
  wire             _GEN_32 = ~icache_resp.valid | ~dcache_resp.valid;
  reg  [1:0]       Register_inst6;
  reg  [2:0]       Register_inst7;
  reg              Register_inst9;
  reg              Register_inst11;
  reg              Register_inst12;
  reg  [31:0]      Register_inst3;
  wire [1:0][31:0] _GEN_33 = {{Register_inst14}, {Register_inst14 + 32'h4}};
  reg              Register_inst13;
  reg  [31:0]      Register_inst4;
  reg  [31:0]      Register_inst2;
  reg  [1:0]       Register_inst8;
  wire             rs2_hazard =
    Register_inst9 & (|(Register_inst0[24:20]))
    & Register_inst0[24:20] == Register_inst2[11:7] & Register_inst8 == 2'h0;
  wire [1:0][31:0] _GEN_34 = {{Register_inst4}, {_RegFile_inst0_rdata2}};
  wire             is_nop =
    Register_inst13 | ctrl_inst_kill | _BrCondArea_inst0_taken | _CSRGen_inst0_expt;
  wire [31:0]      _GEN_35 = dcache_resp.data.data >> {27'h0, Register_inst4[1:0], 3'h0};
  wire [1:0][31:0] _GEN_36 =
    {{{{17{_GEN_35[15]}}, _GEN_35[14:0]}}, {dcache_resp.data.data}};
  wire [1:0][31:0] _GEN_37 =
    {{{16'h0, _GEN_35[15:0]}}, {_GEN_36[Register_inst7 == 3'h2]}};
  wire [1:0][31:0] _GEN_38 =
    {{{{25{_GEN_35[7]}}, _GEN_35[6:0]}}, {_GEN_37[Register_inst7 == 3'h4]}};
  wire [1:0][31:0] _GEN_39 = {{{24'h0, _GEN_35[7:0]}}, {_GEN_38[Register_inst7 == 3'h3]}};
  wire [1:0][31:0] _GEN_40 = {{_GEN_39[Register_inst7 == 3'h5]}, {Register_inst4}};
  wire [1:0][31:0] _GEN_41 =
    {{Register_inst3 + 32'h4}, {_GEN_40[Register_inst8 == 2'h1]}};
  wire [1:0][31:0] _GEN_42 = {{_CSRGen_inst0_O}, {_GEN_41[Register_inst8 == 2'h2]}};
  wire             rs1_hazard =
    Register_inst9 & (|(Register_inst0[19:15]))
    & Register_inst0[19:15] == Register_inst2[11:7] & Register_inst8 == 2'h0;
  wire [1:0][31:0] _GEN_43 = {{Register_inst4}, {_RegFile_inst0_rdata1}};
  wire [1:0][31:0] _GEN_44 = {{_GEN_43[rs1_hazard]}, {Register_inst1}};
  wire [1:0][31:0] _GEN_45 = {{_GEN_34[rs2_hazard]}, {_ImmGenWire_inst0_O}};
  wire             take_sum = ctrl_pc_sel == 2'h1 | _BrCondArea_inst0_taken;
  wire [1:0][31:0] _GEN_46 =
    {{{_ALUArea_inst0_sum_[31:1], 1'h0}}, {_GEN_33[ctrl_pc_sel == 2'h2]}};
  wire [1:0][31:0] _GEN_47 = {{_CSRGen_inst0_epc}, {_GEN_46[take_sum]}};
  wire [1:0][31:0] _GEN_48 = {{_CSRGen_inst0_evec}, {_GEN_47[&ctrl_pc_sel]}};
  wire [1:0][31:0] _GEN_49 = {{Register_inst14}, {_GEN_48[_CSRGen_inst0_expt]}};
  wire [1:0][31:0] _GEN_50 = {{32'h13}, {icache_resp.data.data}};
  always_ff @(posedge CLK) begin
    if (RESET) begin
      Register_inst2 <= 32'h13;
      Register_inst0 <= 32'h13;
      Register_inst14 <= 32'h1FC;
    end
    else begin
      Register_inst2 <=
        {_GEN,
         _GEN_0,
         _GEN_1,
         _GEN_2,
         _GEN_3,
         _GEN_4,
         _GEN_5,
         _GEN_6,
         _GEN_7,
         _GEN_8,
         _GEN_9,
         _GEN_10,
         _GEN_11,
         _GEN_12,
         _GEN_13,
         _GEN_14,
         _GEN_15,
         _GEN_16,
         _GEN_17,
         _GEN_18,
         _GEN_19,
         _GEN_20,
         _GEN_21,
         _GEN_22,
         _GEN_23,
         _GEN_24,
         _GEN_25,
         _GEN_26,
         _GEN_27,
         _GEN_28,
         _GEN_29,
         _GEN_30};
      if (~_GEN_32)
        Register_inst0 <= _GEN_50[is_nop];
      Register_inst14 <= _GEN_49[_GEN_32];
    end
  end // always_ff @(posedge)
  reg  [31:0]      Register_inst5;
  reg  [1:0]       _GEN_51;
  reg  [2:0]       _GEN_52;
  reg              _GEN_53;
  reg  [2:0]       _GEN_54;
  reg              _GEN_55;
  reg              _GEN_56;
  reg  [31:0]      _GEN_57;
  reg  [31:0]      _GEN_58;
  reg  [31:0]      _GEN_59;
  reg  [1:0]       _GEN_60;
  wire [1:0][31:0] _GEN_61 = {{_ImmGenWire_inst0_O}, {_GEN_43[rs1_hazard]}};
  always_comb begin
    _GEN_51 = Register_inst6;
    _GEN_52 = Register_inst7;
    _GEN_53 = Register_inst9;
    _GEN_54 = Register_inst10;
    _GEN_55 = Register_inst11;
    _GEN_56 = Register_inst12;
    _GEN_57 = Register_inst3;
    _GEN_30 = Register_inst2[0];
    _GEN_29 = Register_inst2[1];
    _GEN_28 = Register_inst2[2];
    _GEN_27 = Register_inst2[3];
    _GEN_26 = Register_inst2[4];
    _GEN_25 = Register_inst2[5];
    _GEN_24 = Register_inst2[6];
    _GEN_23 = Register_inst2[7];
    _GEN_22 = Register_inst2[8];
    _GEN_21 = Register_inst2[9];
    _GEN_20 = Register_inst2[10];
    _GEN_19 = Register_inst2[11];
    _GEN_18 = Register_inst2[12];
    _GEN_17 = Register_inst2[13];
    _GEN_16 = Register_inst2[14];
    _GEN_15 = Register_inst2[15];
    _GEN_14 = Register_inst2[16];
    _GEN_13 = Register_inst2[17];
    _GEN_12 = Register_inst2[18];
    _GEN_11 = Register_inst2[19];
    _GEN_10 = Register_inst2[20];
    _GEN_9 = Register_inst2[21];
    _GEN_8 = Register_inst2[22];
    _GEN_7 = Register_inst2[23];
    _GEN_6 = Register_inst2[24];
    _GEN_5 = Register_inst2[25];
    _GEN_4 = Register_inst2[26];
    _GEN_3 = Register_inst2[27];
    _GEN_2 = Register_inst2[28];
    _GEN_1 = Register_inst2[29];
    _GEN_0 = Register_inst2[30];
    _GEN = Register_inst2[31];
    _GEN_58 = Register_inst4;
    _GEN_59 = Register_inst5;
    _GEN_60 = Register_inst8;
    if (RESET | ~_GEN_32 & _CSRGen_inst0_expt) begin
      _GEN_51 = 2'h0;
      _GEN_52 = 3'h0;
      _GEN_53 = 1'h0;
      _GEN_54 = 3'h0;
      _GEN_55 = 1'h0;
      _GEN_56 = 1'h0;
    end
    else if (~_GEN_32 & ~_CSRGen_inst0_expt) begin
      _GEN_57 = Register_inst1;
      _GEN_30 = Register_inst0[0];
      _GEN_29 = Register_inst0[1];
      _GEN_28 = Register_inst0[2];
      _GEN_27 = Register_inst0[3];
      _GEN_26 = Register_inst0[4];
      _GEN_25 = Register_inst0[5];
      _GEN_24 = Register_inst0[6];
      _GEN_23 = Register_inst0[7];
      _GEN_22 = Register_inst0[8];
      _GEN_21 = Register_inst0[9];
      _GEN_20 = Register_inst0[10];
      _GEN_19 = Register_inst0[11];
      _GEN_18 = Register_inst0[12];
      _GEN_17 = Register_inst0[13];
      _GEN_16 = Register_inst0[14];
      _GEN_15 = Register_inst0[15];
      _GEN_14 = Register_inst0[16];
      _GEN_13 = Register_inst0[17];
      _GEN_12 = Register_inst0[18];
      _GEN_11 = Register_inst0[19];
      _GEN_10 = Register_inst0[20];
      _GEN_9 = Register_inst0[21];
      _GEN_8 = Register_inst0[22];
      _GEN_7 = Register_inst0[23];
      _GEN_6 = Register_inst0[24];
      _GEN_5 = Register_inst0[25];
      _GEN_4 = Register_inst0[26];
      _GEN_3 = Register_inst0[27];
      _GEN_2 = Register_inst0[28];
      _GEN_1 = Register_inst0[29];
      _GEN_0 = Register_inst0[30];
      _GEN = Register_inst0[31];
      _GEN_58 = _ALUArea_inst0_O;
      _GEN_59 = _GEN_61[ctrl_imm_sel == 3'h6];
      _GEN_51 = ctrl_st_type;
      _GEN_52 = ctrl_ld_type;
      _GEN_60 = ctrl_wb_sel;
      _GEN_53 = ctrl_wb_en;
      _GEN_54 = ctrl_csr_cmd;
      _GEN_55 = ctrl_illegal;
      _GEN_56 = ctrl_pc_sel == 2'h1;
    end
  end // always_comb
  always_ff @(posedge CLK) begin
    Register_inst6 <= _GEN_51;
    Register_inst7 <= _GEN_52;
    Register_inst9 <= _GEN_53;
    Register_inst11 <= _GEN_55;
    Register_inst12 <= _GEN_56;
    Register_inst3 <= _GEN_57;
    Register_inst13 <= RESET;
    Register_inst4 <= _GEN_58;
    Register_inst8 <= _GEN_60;
    if (~_GEN_32)
      Register_inst1 <= Register_inst14;
    Register_inst5 <= _GEN_59;
    Register_inst10 <= _GEN_54;
  end // always_ff @(posedge)
  initial begin
    Register_inst6 = 2'h0;
    Register_inst7 = 3'h0;
    Register_inst9 = 1'h0;
    Register_inst11 = 1'h0;
    Register_inst12 = 1'h0;
    Register_inst3 = 32'h0;
    Register_inst13 = 1'h0;
    Register_inst4 = 32'h0;
    Register_inst2 = 32'h13;
    Register_inst8 = 2'h0;
    Register_inst0 = 32'h13;
    Register_inst14 = 32'h1FC;
    Register_inst1 = 32'h0;
    Register_inst5 = 32'h0;
    Register_inst10 = 3'h0;
  end // initial
  wire struct packed {logic [31:0] addr; logic [31:0] data; logic [3:0] mask; } _GEN_62;
  assign _GEN_62.addr = _GEN_49[_GEN_32];
  assign _GEN_62.data = 32'h0;
  assign _GEN_62.mask = 4'h0;
  wire
    struct packed {logic valid; struct packed {logic [31:0] addr; logic [31:0] data; logic [3:0] mask; } data; }
    _GEN_63;
  assign _GEN_63.valid = ~_GEN_32;
  assign _GEN_63.data = _GEN_62;
  wire [1:0][31:0] _GEN_64 = {{Register_inst4}, {_ALUArea_inst0_sum_}};
  wire [1:0][1:0]  _GEN_65 = {{Register_inst6}, {ctrl_st_type}};
  wire [1:0][3:0]  _GEN_66 =
    {{4'h3 << _ALUArea_inst0_sum_[1:0]}, {_GEN_31[_GEN_65[_GEN_32] == 2'h1]}};
  wire [1:0][3:0]  _GEN_67 =
    {{4'h1 << _ALUArea_inst0_sum_[1:0]}, {_GEN_66[_GEN_65[_GEN_32] == 2'h2]}};
  wire struct packed {logic [31:0] addr; logic [31:0] data; logic [3:0] mask; } _GEN_68;
  assign _GEN_68.addr = {_GEN_64[_GEN_32][31:2], 2'h0};
  assign _GEN_68.data = _GEN_34[rs2_hazard] << {27'h0, _ALUArea_inst0_sum_[1:0], 3'h0};
  assign _GEN_68.mask = _GEN_67[&_GEN_65[_GEN_32]];
  wire
    struct packed {logic valid; struct packed {logic [31:0] addr; logic [31:0] data; logic [3:0] mask; } data; }
    _GEN_69;
  assign _GEN_69.valid = ~_GEN_32 & ((|ctrl_st_type) | (|ctrl_ld_type));
  assign _GEN_69.data = _GEN_68;
  BrCondArea BrCondArea_inst0 (
    .rs1     (_GEN_43[rs1_hazard]),
    .rs2     (_GEN_34[rs2_hazard]),
    .br_type (ctrl_br_type),
    .taken   (_BrCondArea_inst0_taken)
  );
  RegFile RegFile_inst0 (
    .raddr1 (Register_inst0[19:15]),
    .raddr2 (Register_inst0[24:20]),
    .wen    (Register_inst9 & ~_GEN_32 & ~_CSRGen_inst0_expt),
    .waddr  (Register_inst2[11:7]),
    .wdata  (_GEN_42[&Register_inst8]),
    .CLK    (CLK),
    .RESET  (RESET),
    .rdata1 (_RegFile_inst0_rdata1),
    .rdata2 (_RegFile_inst0_rdata2)
  );
  ImmGenWire ImmGenWire_inst0 (
    .inst (Register_inst0),
    .sel  (ctrl_imm_sel),
    .O    (_ImmGenWire_inst0_O)
  );
  ALUArea ALUArea_inst0 (
    .A    (_GEN_44[ctrl_A_sel]),
    .B    (_GEN_45[ctrl_B_sel]),
    .op   (ctrl_alu_op),
    .O    (_ALUArea_inst0_O),
    .sum_ (_ALUArea_inst0_sum_)
  );
  CSRGen CSRGen_inst0 (
    .stall         (_GEN_32),
    .cmd           (Register_inst10),
    .I             (Register_inst5),
    .pc            (Register_inst3),
    .addr          (Register_inst4),
    .inst          (Register_inst2),
    .illegal       (Register_inst11),
    .st_type       (Register_inst6),
    .ld_type       (Register_inst7),
    .pc_check      (Register_inst12),
    .host_fromhost (host_fromhost),
    .CLK           (CLK),
    .RESET         (RESET),
    .O             (_CSRGen_inst0_O),
    .expt          (_CSRGen_inst0_expt),
    .evec          (_CSRGen_inst0_evec),
    .epc           (_CSRGen_inst0_epc),
    .host_tohost   (host_tohost)
  );
  assign icache_abort = 1'h0;
  assign icache_req = _GEN_63;
  assign dcache_abort = _CSRGen_inst0_expt;
  assign dcache_req = _GEN_69;
  assign ctrl_inst = Register_inst0;
endmodule

module Control(
  input  [31:0] inst,
  output [1:0]  pc_sel,
  output        inst_kill,
                A_sel,
                B_sel,
  output [2:0]  imm_sel,
  output [3:0]  alu_op,
  output [2:0]  br_type,
  output [1:0]  st_type,
  output [2:0]  ld_type,
  output [1:0]  wb_sel,
  output        wb_en,
  output [2:0]  csr_cmd,
  output        illegal
);

  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN;
  assign _GEN._0 = 2'h0;
  assign _GEN._1 = 1'h0;
  assign _GEN._2 = 1'h0;
  assign _GEN._3 = 3'h0;
  assign _GEN._4 = 4'hF;
  assign _GEN._5 = 3'h0;
  assign _GEN._6 = 1'h0;
  assign _GEN._7 = 2'h0;
  assign _GEN._8 = 3'h0;
  assign _GEN._9 = 2'h0;
  assign _GEN._10 = 1'h0;
  assign _GEN._11 = 3'h0;
  assign _GEN._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_0;
  assign _GEN_0._0 = 2'h3;
  assign _GEN_0._1 = 1'h0;
  assign _GEN_0._2 = 1'h0;
  assign _GEN_0._3 = 3'h0;
  assign _GEN_0._4 = 4'hF;
  assign _GEN_0._5 = 3'h0;
  assign _GEN_0._6 = 1'h1;
  assign _GEN_0._7 = 2'h0;
  assign _GEN_0._8 = 3'h0;
  assign _GEN_0._9 = 2'h3;
  assign _GEN_0._10 = 1'h0;
  assign _GEN_0._11 = 3'h4;
  assign _GEN_0._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_1;
  assign _GEN_1._0 = 2'h0;
  assign _GEN_1._1 = 1'h0;
  assign _GEN_1._2 = 1'h0;
  assign _GEN_1._3 = 3'h0;
  assign _GEN_1._4 = 4'hF;
  assign _GEN_1._5 = 3'h0;
  assign _GEN_1._6 = 1'h0;
  assign _GEN_1._7 = 2'h0;
  assign _GEN_1._8 = 3'h0;
  assign _GEN_1._9 = 2'h3;
  assign _GEN_1._10 = 1'h0;
  assign _GEN_1._11 = 3'h4;
  assign _GEN_1._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_2;
  assign _GEN_2._0 = 2'h2;
  assign _GEN_2._1 = 1'h0;
  assign _GEN_2._2 = 1'h0;
  assign _GEN_2._3 = 3'h6;
  assign _GEN_2._4 = 4'hF;
  assign _GEN_2._5 = 3'h0;
  assign _GEN_2._6 = 1'h1;
  assign _GEN_2._7 = 2'h0;
  assign _GEN_2._8 = 3'h0;
  assign _GEN_2._9 = 2'h3;
  assign _GEN_2._10 = 1'h1;
  assign _GEN_2._11 = 3'h3;
  assign _GEN_2._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_3;
  assign _GEN_3._0 = 2'h2;
  assign _GEN_3._1 = 1'h0;
  assign _GEN_3._2 = 1'h0;
  assign _GEN_3._3 = 3'h6;
  assign _GEN_3._4 = 4'hF;
  assign _GEN_3._5 = 3'h0;
  assign _GEN_3._6 = 1'h1;
  assign _GEN_3._7 = 2'h0;
  assign _GEN_3._8 = 3'h0;
  assign _GEN_3._9 = 2'h3;
  assign _GEN_3._10 = 1'h1;
  assign _GEN_3._11 = 3'h2;
  assign _GEN_3._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_4;
  assign _GEN_4._0 = 2'h2;
  assign _GEN_4._1 = 1'h0;
  assign _GEN_4._2 = 1'h0;
  assign _GEN_4._3 = 3'h6;
  assign _GEN_4._4 = 4'hF;
  assign _GEN_4._5 = 3'h0;
  assign _GEN_4._6 = 1'h1;
  assign _GEN_4._7 = 2'h0;
  assign _GEN_4._8 = 3'h0;
  assign _GEN_4._9 = 2'h3;
  assign _GEN_4._10 = 1'h1;
  assign _GEN_4._11 = 3'h1;
  assign _GEN_4._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_5;
  assign _GEN_5._0 = 2'h2;
  assign _GEN_5._1 = 1'h1;
  assign _GEN_5._2 = 1'h0;
  assign _GEN_5._3 = 3'h0;
  assign _GEN_5._4 = 4'hA;
  assign _GEN_5._5 = 3'h0;
  assign _GEN_5._6 = 1'h1;
  assign _GEN_5._7 = 2'h0;
  assign _GEN_5._8 = 3'h0;
  assign _GEN_5._9 = 2'h3;
  assign _GEN_5._10 = 1'h1;
  assign _GEN_5._11 = 3'h3;
  assign _GEN_5._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_6;
  assign _GEN_6._0 = 2'h2;
  assign _GEN_6._1 = 1'h1;
  assign _GEN_6._2 = 1'h0;
  assign _GEN_6._3 = 3'h0;
  assign _GEN_6._4 = 4'hA;
  assign _GEN_6._5 = 3'h0;
  assign _GEN_6._6 = 1'h1;
  assign _GEN_6._7 = 2'h0;
  assign _GEN_6._8 = 3'h0;
  assign _GEN_6._9 = 2'h3;
  assign _GEN_6._10 = 1'h1;
  assign _GEN_6._11 = 3'h2;
  assign _GEN_6._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_7;
  assign _GEN_7._0 = 2'h2;
  assign _GEN_7._1 = 1'h1;
  assign _GEN_7._2 = 1'h0;
  assign _GEN_7._3 = 3'h0;
  assign _GEN_7._4 = 4'hA;
  assign _GEN_7._5 = 3'h0;
  assign _GEN_7._6 = 1'h1;
  assign _GEN_7._7 = 2'h0;
  assign _GEN_7._8 = 3'h0;
  assign _GEN_7._9 = 2'h3;
  assign _GEN_7._10 = 1'h1;
  assign _GEN_7._11 = 3'h1;
  assign _GEN_7._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_8;
  assign _GEN_8._0 = 2'h2;
  assign _GEN_8._1 = 1'h0;
  assign _GEN_8._2 = 1'h0;
  assign _GEN_8._3 = 3'h0;
  assign _GEN_8._4 = 4'hF;
  assign _GEN_8._5 = 3'h0;
  assign _GEN_8._6 = 1'h1;
  assign _GEN_8._7 = 2'h0;
  assign _GEN_8._8 = 3'h0;
  assign _GEN_8._9 = 2'h0;
  assign _GEN_8._10 = 1'h0;
  assign _GEN_8._11 = 3'h0;
  assign _GEN_8._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_9;
  assign _GEN_9._0 = 2'h0;
  assign _GEN_9._1 = 1'h1;
  assign _GEN_9._2 = 1'h1;
  assign _GEN_9._3 = 3'h0;
  assign _GEN_9._4 = 4'h2;
  assign _GEN_9._5 = 3'h0;
  assign _GEN_9._6 = 1'h0;
  assign _GEN_9._7 = 2'h0;
  assign _GEN_9._8 = 3'h0;
  assign _GEN_9._9 = 2'h0;
  assign _GEN_9._10 = 1'h1;
  assign _GEN_9._11 = 3'h0;
  assign _GEN_9._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_10;
  assign _GEN_10._0 = 2'h0;
  assign _GEN_10._1 = 1'h1;
  assign _GEN_10._2 = 1'h1;
  assign _GEN_10._3 = 3'h0;
  assign _GEN_10._4 = 4'h3;
  assign _GEN_10._5 = 3'h0;
  assign _GEN_10._6 = 1'h0;
  assign _GEN_10._7 = 2'h0;
  assign _GEN_10._8 = 3'h0;
  assign _GEN_10._9 = 2'h0;
  assign _GEN_10._10 = 1'h1;
  assign _GEN_10._11 = 3'h0;
  assign _GEN_10._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_11;
  assign _GEN_11._0 = 2'h0;
  assign _GEN_11._1 = 1'h1;
  assign _GEN_11._2 = 1'h1;
  assign _GEN_11._3 = 3'h0;
  assign _GEN_11._4 = 4'h9;
  assign _GEN_11._5 = 3'h0;
  assign _GEN_11._6 = 1'h0;
  assign _GEN_11._7 = 2'h0;
  assign _GEN_11._8 = 3'h0;
  assign _GEN_11._9 = 2'h0;
  assign _GEN_11._10 = 1'h1;
  assign _GEN_11._11 = 3'h0;
  assign _GEN_11._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_12;
  assign _GEN_12._0 = 2'h0;
  assign _GEN_12._1 = 1'h1;
  assign _GEN_12._2 = 1'h1;
  assign _GEN_12._3 = 3'h0;
  assign _GEN_12._4 = 4'h8;
  assign _GEN_12._5 = 3'h0;
  assign _GEN_12._6 = 1'h0;
  assign _GEN_12._7 = 2'h0;
  assign _GEN_12._8 = 3'h0;
  assign _GEN_12._9 = 2'h0;
  assign _GEN_12._10 = 1'h1;
  assign _GEN_12._11 = 3'h0;
  assign _GEN_12._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_13;
  assign _GEN_13._0 = 2'h0;
  assign _GEN_13._1 = 1'h1;
  assign _GEN_13._2 = 1'h1;
  assign _GEN_13._3 = 3'h0;
  assign _GEN_13._4 = 4'h4;
  assign _GEN_13._5 = 3'h0;
  assign _GEN_13._6 = 1'h0;
  assign _GEN_13._7 = 2'h0;
  assign _GEN_13._8 = 3'h0;
  assign _GEN_13._9 = 2'h0;
  assign _GEN_13._10 = 1'h1;
  assign _GEN_13._11 = 3'h0;
  assign _GEN_13._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_14;
  assign _GEN_14._0 = 2'h0;
  assign _GEN_14._1 = 1'h1;
  assign _GEN_14._2 = 1'h1;
  assign _GEN_14._3 = 3'h0;
  assign _GEN_14._4 = 4'h7;
  assign _GEN_14._5 = 3'h0;
  assign _GEN_14._6 = 1'h0;
  assign _GEN_14._7 = 2'h0;
  assign _GEN_14._8 = 3'h0;
  assign _GEN_14._9 = 2'h0;
  assign _GEN_14._10 = 1'h1;
  assign _GEN_14._11 = 3'h0;
  assign _GEN_14._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_15;
  assign _GEN_15._0 = 2'h0;
  assign _GEN_15._1 = 1'h1;
  assign _GEN_15._2 = 1'h1;
  assign _GEN_15._3 = 3'h0;
  assign _GEN_15._4 = 4'h5;
  assign _GEN_15._5 = 3'h0;
  assign _GEN_15._6 = 1'h0;
  assign _GEN_15._7 = 2'h0;
  assign _GEN_15._8 = 3'h0;
  assign _GEN_15._9 = 2'h0;
  assign _GEN_15._10 = 1'h1;
  assign _GEN_15._11 = 3'h0;
  assign _GEN_15._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_16;
  assign _GEN_16._0 = 2'h0;
  assign _GEN_16._1 = 1'h1;
  assign _GEN_16._2 = 1'h1;
  assign _GEN_16._3 = 3'h0;
  assign _GEN_16._4 = 4'h6;
  assign _GEN_16._5 = 3'h0;
  assign _GEN_16._6 = 1'h0;
  assign _GEN_16._7 = 2'h0;
  assign _GEN_16._8 = 3'h0;
  assign _GEN_16._9 = 2'h0;
  assign _GEN_16._10 = 1'h1;
  assign _GEN_16._11 = 3'h0;
  assign _GEN_16._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_17;
  assign _GEN_17._0 = 2'h0;
  assign _GEN_17._1 = 1'h1;
  assign _GEN_17._2 = 1'h1;
  assign _GEN_17._3 = 3'h0;
  assign _GEN_17._4 = 4'h1;
  assign _GEN_17._5 = 3'h0;
  assign _GEN_17._6 = 1'h0;
  assign _GEN_17._7 = 2'h0;
  assign _GEN_17._8 = 3'h0;
  assign _GEN_17._9 = 2'h0;
  assign _GEN_17._10 = 1'h1;
  assign _GEN_17._11 = 3'h0;
  assign _GEN_17._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_18;
  assign _GEN_18._0 = 2'h0;
  assign _GEN_18._1 = 1'h1;
  assign _GEN_18._2 = 1'h1;
  assign _GEN_18._3 = 3'h0;
  assign _GEN_18._4 = 4'h0;
  assign _GEN_18._5 = 3'h0;
  assign _GEN_18._6 = 1'h0;
  assign _GEN_18._7 = 2'h0;
  assign _GEN_18._8 = 3'h0;
  assign _GEN_18._9 = 2'h0;
  assign _GEN_18._10 = 1'h1;
  assign _GEN_18._11 = 3'h0;
  assign _GEN_18._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_19;
  assign _GEN_19._0 = 2'h0;
  assign _GEN_19._1 = 1'h1;
  assign _GEN_19._2 = 1'h0;
  assign _GEN_19._3 = 3'h1;
  assign _GEN_19._4 = 4'h9;
  assign _GEN_19._5 = 3'h0;
  assign _GEN_19._6 = 1'h0;
  assign _GEN_19._7 = 2'h0;
  assign _GEN_19._8 = 3'h0;
  assign _GEN_19._9 = 2'h0;
  assign _GEN_19._10 = 1'h1;
  assign _GEN_19._11 = 3'h0;
  assign _GEN_19._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_20;
  assign _GEN_20._0 = 2'h0;
  assign _GEN_20._1 = 1'h1;
  assign _GEN_20._2 = 1'h0;
  assign _GEN_20._3 = 3'h1;
  assign _GEN_20._4 = 4'h8;
  assign _GEN_20._5 = 3'h0;
  assign _GEN_20._6 = 1'h0;
  assign _GEN_20._7 = 2'h0;
  assign _GEN_20._8 = 3'h0;
  assign _GEN_20._9 = 2'h0;
  assign _GEN_20._10 = 1'h1;
  assign _GEN_20._11 = 3'h0;
  assign _GEN_20._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_21;
  assign _GEN_21._0 = 2'h0;
  assign _GEN_21._1 = 1'h1;
  assign _GEN_21._2 = 1'h0;
  assign _GEN_21._3 = 3'h1;
  assign _GEN_21._4 = 4'h6;
  assign _GEN_21._5 = 3'h0;
  assign _GEN_21._6 = 1'h0;
  assign _GEN_21._7 = 2'h0;
  assign _GEN_21._8 = 3'h0;
  assign _GEN_21._9 = 2'h0;
  assign _GEN_21._10 = 1'h1;
  assign _GEN_21._11 = 3'h0;
  assign _GEN_21._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_22;
  assign _GEN_22._0 = 2'h0;
  assign _GEN_22._1 = 1'h1;
  assign _GEN_22._2 = 1'h0;
  assign _GEN_22._3 = 3'h1;
  assign _GEN_22._4 = 4'h2;
  assign _GEN_22._5 = 3'h0;
  assign _GEN_22._6 = 1'h0;
  assign _GEN_22._7 = 2'h0;
  assign _GEN_22._8 = 3'h0;
  assign _GEN_22._9 = 2'h0;
  assign _GEN_22._10 = 1'h1;
  assign _GEN_22._11 = 3'h0;
  assign _GEN_22._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_23;
  assign _GEN_23._0 = 2'h0;
  assign _GEN_23._1 = 1'h1;
  assign _GEN_23._2 = 1'h0;
  assign _GEN_23._3 = 3'h1;
  assign _GEN_23._4 = 4'h3;
  assign _GEN_23._5 = 3'h0;
  assign _GEN_23._6 = 1'h0;
  assign _GEN_23._7 = 2'h0;
  assign _GEN_23._8 = 3'h0;
  assign _GEN_23._9 = 2'h0;
  assign _GEN_23._10 = 1'h1;
  assign _GEN_23._11 = 3'h0;
  assign _GEN_23._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_24;
  assign _GEN_24._0 = 2'h0;
  assign _GEN_24._1 = 1'h1;
  assign _GEN_24._2 = 1'h0;
  assign _GEN_24._3 = 3'h1;
  assign _GEN_24._4 = 4'h4;
  assign _GEN_24._5 = 3'h0;
  assign _GEN_24._6 = 1'h0;
  assign _GEN_24._7 = 2'h0;
  assign _GEN_24._8 = 3'h0;
  assign _GEN_24._9 = 2'h0;
  assign _GEN_24._10 = 1'h1;
  assign _GEN_24._11 = 3'h0;
  assign _GEN_24._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_25;
  assign _GEN_25._0 = 2'h0;
  assign _GEN_25._1 = 1'h1;
  assign _GEN_25._2 = 1'h0;
  assign _GEN_25._3 = 3'h1;
  assign _GEN_25._4 = 4'h7;
  assign _GEN_25._5 = 3'h0;
  assign _GEN_25._6 = 1'h0;
  assign _GEN_25._7 = 2'h0;
  assign _GEN_25._8 = 3'h0;
  assign _GEN_25._9 = 2'h0;
  assign _GEN_25._10 = 1'h1;
  assign _GEN_25._11 = 3'h0;
  assign _GEN_25._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_26;
  assign _GEN_26._0 = 2'h0;
  assign _GEN_26._1 = 1'h1;
  assign _GEN_26._2 = 1'h0;
  assign _GEN_26._3 = 3'h1;
  assign _GEN_26._4 = 4'h5;
  assign _GEN_26._5 = 3'h0;
  assign _GEN_26._6 = 1'h0;
  assign _GEN_26._7 = 2'h0;
  assign _GEN_26._8 = 3'h0;
  assign _GEN_26._9 = 2'h0;
  assign _GEN_26._10 = 1'h1;
  assign _GEN_26._11 = 3'h0;
  assign _GEN_26._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_27;
  assign _GEN_27._0 = 2'h0;
  assign _GEN_27._1 = 1'h1;
  assign _GEN_27._2 = 1'h0;
  assign _GEN_27._3 = 3'h1;
  assign _GEN_27._4 = 4'h0;
  assign _GEN_27._5 = 3'h0;
  assign _GEN_27._6 = 1'h0;
  assign _GEN_27._7 = 2'h0;
  assign _GEN_27._8 = 3'h0;
  assign _GEN_27._9 = 2'h0;
  assign _GEN_27._10 = 1'h1;
  assign _GEN_27._11 = 3'h0;
  assign _GEN_27._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_28;
  assign _GEN_28._0 = 2'h0;
  assign _GEN_28._1 = 1'h1;
  assign _GEN_28._2 = 1'h0;
  assign _GEN_28._3 = 3'h2;
  assign _GEN_28._4 = 4'h0;
  assign _GEN_28._5 = 3'h0;
  assign _GEN_28._6 = 1'h0;
  assign _GEN_28._7 = 2'h1;
  assign _GEN_28._8 = 3'h0;
  assign _GEN_28._9 = 2'h0;
  assign _GEN_28._10 = 1'h0;
  assign _GEN_28._11 = 3'h0;
  assign _GEN_28._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_29;
  assign _GEN_29._0 = 2'h0;
  assign _GEN_29._1 = 1'h1;
  assign _GEN_29._2 = 1'h0;
  assign _GEN_29._3 = 3'h2;
  assign _GEN_29._4 = 4'h0;
  assign _GEN_29._5 = 3'h0;
  assign _GEN_29._6 = 1'h0;
  assign _GEN_29._7 = 2'h2;
  assign _GEN_29._8 = 3'h0;
  assign _GEN_29._9 = 2'h0;
  assign _GEN_29._10 = 1'h0;
  assign _GEN_29._11 = 3'h0;
  assign _GEN_29._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_30;
  assign _GEN_30._0 = 2'h0;
  assign _GEN_30._1 = 1'h1;
  assign _GEN_30._2 = 1'h0;
  assign _GEN_30._3 = 3'h2;
  assign _GEN_30._4 = 4'h0;
  assign _GEN_30._5 = 3'h0;
  assign _GEN_30._6 = 1'h0;
  assign _GEN_30._7 = 2'h3;
  assign _GEN_30._8 = 3'h0;
  assign _GEN_30._9 = 2'h0;
  assign _GEN_30._10 = 1'h0;
  assign _GEN_30._11 = 3'h0;
  assign _GEN_30._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_31;
  assign _GEN_31._0 = 2'h2;
  assign _GEN_31._1 = 1'h1;
  assign _GEN_31._2 = 1'h0;
  assign _GEN_31._3 = 3'h1;
  assign _GEN_31._4 = 4'h0;
  assign _GEN_31._5 = 3'h0;
  assign _GEN_31._6 = 1'h1;
  assign _GEN_31._7 = 2'h0;
  assign _GEN_31._8 = 3'h4;
  assign _GEN_31._9 = 2'h1;
  assign _GEN_31._10 = 1'h1;
  assign _GEN_31._11 = 3'h0;
  assign _GEN_31._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_32;
  assign _GEN_32._0 = 2'h2;
  assign _GEN_32._1 = 1'h1;
  assign _GEN_32._2 = 1'h0;
  assign _GEN_32._3 = 3'h1;
  assign _GEN_32._4 = 4'h0;
  assign _GEN_32._5 = 3'h0;
  assign _GEN_32._6 = 1'h1;
  assign _GEN_32._7 = 2'h0;
  assign _GEN_32._8 = 3'h5;
  assign _GEN_32._9 = 2'h1;
  assign _GEN_32._10 = 1'h1;
  assign _GEN_32._11 = 3'h0;
  assign _GEN_32._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_33;
  assign _GEN_33._0 = 2'h2;
  assign _GEN_33._1 = 1'h1;
  assign _GEN_33._2 = 1'h0;
  assign _GEN_33._3 = 3'h1;
  assign _GEN_33._4 = 4'h0;
  assign _GEN_33._5 = 3'h0;
  assign _GEN_33._6 = 1'h1;
  assign _GEN_33._7 = 2'h0;
  assign _GEN_33._8 = 3'h1;
  assign _GEN_33._9 = 2'h1;
  assign _GEN_33._10 = 1'h1;
  assign _GEN_33._11 = 3'h0;
  assign _GEN_33._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_34;
  assign _GEN_34._0 = 2'h2;
  assign _GEN_34._1 = 1'h1;
  assign _GEN_34._2 = 1'h0;
  assign _GEN_34._3 = 3'h1;
  assign _GEN_34._4 = 4'h0;
  assign _GEN_34._5 = 3'h0;
  assign _GEN_34._6 = 1'h1;
  assign _GEN_34._7 = 2'h0;
  assign _GEN_34._8 = 3'h2;
  assign _GEN_34._9 = 2'h1;
  assign _GEN_34._10 = 1'h1;
  assign _GEN_34._11 = 3'h0;
  assign _GEN_34._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_35;
  assign _GEN_35._0 = 2'h2;
  assign _GEN_35._1 = 1'h1;
  assign _GEN_35._2 = 1'h0;
  assign _GEN_35._3 = 3'h1;
  assign _GEN_35._4 = 4'h0;
  assign _GEN_35._5 = 3'h0;
  assign _GEN_35._6 = 1'h1;
  assign _GEN_35._7 = 2'h0;
  assign _GEN_35._8 = 3'h3;
  assign _GEN_35._9 = 2'h1;
  assign _GEN_35._10 = 1'h1;
  assign _GEN_35._11 = 3'h0;
  assign _GEN_35._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_36;
  assign _GEN_36._0 = 2'h0;
  assign _GEN_36._1 = 1'h0;
  assign _GEN_36._2 = 1'h0;
  assign _GEN_36._3 = 3'h5;
  assign _GEN_36._4 = 4'h0;
  assign _GEN_36._5 = 3'h4;
  assign _GEN_36._6 = 1'h0;
  assign _GEN_36._7 = 2'h0;
  assign _GEN_36._8 = 3'h0;
  assign _GEN_36._9 = 2'h0;
  assign _GEN_36._10 = 1'h0;
  assign _GEN_36._11 = 3'h0;
  assign _GEN_36._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_37;
  assign _GEN_37._0 = 2'h0;
  assign _GEN_37._1 = 1'h0;
  assign _GEN_37._2 = 1'h0;
  assign _GEN_37._3 = 3'h5;
  assign _GEN_37._4 = 4'h0;
  assign _GEN_37._5 = 3'h1;
  assign _GEN_37._6 = 1'h0;
  assign _GEN_37._7 = 2'h0;
  assign _GEN_37._8 = 3'h0;
  assign _GEN_37._9 = 2'h0;
  assign _GEN_37._10 = 1'h0;
  assign _GEN_37._11 = 3'h0;
  assign _GEN_37._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_38;
  assign _GEN_38._0 = 2'h0;
  assign _GEN_38._1 = 1'h0;
  assign _GEN_38._2 = 1'h0;
  assign _GEN_38._3 = 3'h5;
  assign _GEN_38._4 = 4'h0;
  assign _GEN_38._5 = 3'h5;
  assign _GEN_38._6 = 1'h0;
  assign _GEN_38._7 = 2'h0;
  assign _GEN_38._8 = 3'h0;
  assign _GEN_38._9 = 2'h0;
  assign _GEN_38._10 = 1'h0;
  assign _GEN_38._11 = 3'h0;
  assign _GEN_38._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_39;
  assign _GEN_39._0 = 2'h0;
  assign _GEN_39._1 = 1'h0;
  assign _GEN_39._2 = 1'h0;
  assign _GEN_39._3 = 3'h5;
  assign _GEN_39._4 = 4'h0;
  assign _GEN_39._5 = 3'h2;
  assign _GEN_39._6 = 1'h0;
  assign _GEN_39._7 = 2'h0;
  assign _GEN_39._8 = 3'h0;
  assign _GEN_39._9 = 2'h0;
  assign _GEN_39._10 = 1'h0;
  assign _GEN_39._11 = 3'h0;
  assign _GEN_39._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_40;
  assign _GEN_40._0 = 2'h0;
  assign _GEN_40._1 = 1'h0;
  assign _GEN_40._2 = 1'h0;
  assign _GEN_40._3 = 3'h5;
  assign _GEN_40._4 = 4'h0;
  assign _GEN_40._5 = 3'h6;
  assign _GEN_40._6 = 1'h0;
  assign _GEN_40._7 = 2'h0;
  assign _GEN_40._8 = 3'h0;
  assign _GEN_40._9 = 2'h0;
  assign _GEN_40._10 = 1'h0;
  assign _GEN_40._11 = 3'h0;
  assign _GEN_40._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_41;
  assign _GEN_41._0 = 2'h0;
  assign _GEN_41._1 = 1'h0;
  assign _GEN_41._2 = 1'h0;
  assign _GEN_41._3 = 3'h5;
  assign _GEN_41._4 = 4'h0;
  assign _GEN_41._5 = 3'h3;
  assign _GEN_41._6 = 1'h0;
  assign _GEN_41._7 = 2'h0;
  assign _GEN_41._8 = 3'h0;
  assign _GEN_41._9 = 2'h0;
  assign _GEN_41._10 = 1'h0;
  assign _GEN_41._11 = 3'h0;
  assign _GEN_41._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_42;
  assign _GEN_42._0 = 2'h1;
  assign _GEN_42._1 = 1'h1;
  assign _GEN_42._2 = 1'h0;
  assign _GEN_42._3 = 3'h1;
  assign _GEN_42._4 = 4'h0;
  assign _GEN_42._5 = 3'h0;
  assign _GEN_42._6 = 1'h1;
  assign _GEN_42._7 = 2'h0;
  assign _GEN_42._8 = 3'h0;
  assign _GEN_42._9 = 2'h2;
  assign _GEN_42._10 = 1'h1;
  assign _GEN_42._11 = 3'h0;
  assign _GEN_42._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_43;
  assign _GEN_43._0 = 2'h1;
  assign _GEN_43._1 = 1'h0;
  assign _GEN_43._2 = 1'h0;
  assign _GEN_43._3 = 3'h4;
  assign _GEN_43._4 = 4'h0;
  assign _GEN_43._5 = 3'h0;
  assign _GEN_43._6 = 1'h1;
  assign _GEN_43._7 = 2'h0;
  assign _GEN_43._8 = 3'h0;
  assign _GEN_43._9 = 2'h2;
  assign _GEN_43._10 = 1'h1;
  assign _GEN_43._11 = 3'h0;
  assign _GEN_43._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_44;
  assign _GEN_44._0 = 2'h0;
  assign _GEN_44._1 = 1'h0;
  assign _GEN_44._2 = 1'h0;
  assign _GEN_44._3 = 3'h3;
  assign _GEN_44._4 = 4'h0;
  assign _GEN_44._5 = 3'h0;
  assign _GEN_44._6 = 1'h0;
  assign _GEN_44._7 = 2'h0;
  assign _GEN_44._8 = 3'h0;
  assign _GEN_44._9 = 2'h0;
  assign _GEN_44._10 = 1'h1;
  assign _GEN_44._11 = 3'h0;
  assign _GEN_44._12 = 1'h0;
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_45 =
    {'{_0: 2'h0,
       _1: 1'h0,
       _2: 1'h0,
       _3: 3'h3,
       _4: 4'hB,
       _5: 3'h0,
       _6: 1'h0,
       _7: 2'h0,
       _8: 3'h0,
       _9: 2'h0,
       _10: 1'h1,
       _11: 3'h0,
       _12: 1'h0},
     '{_0: 2'h0,
       _1: 1'h0,
       _2: 1'h0,
       _3: 3'h0,
       _4: 4'hF,
       _5: 3'h0,
       _6: 1'h0,
       _7: 2'h0,
       _8: 3'h0,
       _9: 2'h0,
       _10: 1'h0,
       _11: 3'h0,
       _12: 1'h1}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_46 = {{_GEN_44}, {_GEN_45[inst[6:0] == 7'h37]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_47 = {{_GEN_43}, {_GEN_46[inst[6:0] == 7'h17]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_48 = {{_GEN_42}, {_GEN_47[inst[6:0] == 7'h6F]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_49 = {{_GEN_41}, {_GEN_48[{inst[14:12], inst[6:0]} == 10'h67]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_50 = {{_GEN_40}, {_GEN_49[{inst[14:12], inst[6:0]} == 10'h63]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_51 = {{_GEN_39}, {_GEN_50[{inst[14:12], inst[6:0]} == 10'hE3]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_52 = {{_GEN_38}, {_GEN_51[{inst[14:12], inst[6:0]} == 10'h263]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_53 = {{_GEN_37}, {_GEN_52[{inst[14:12], inst[6:0]} == 10'h2E3]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_54 = {{_GEN_36}, {_GEN_53[{inst[14:12], inst[6:0]} == 10'h363]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_55 = {{_GEN_35}, {_GEN_54[{inst[14:12], inst[6:0]} == 10'h3E3]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_56 = {{_GEN_34}, {_GEN_55[{inst[14:12], inst[6:0]} == 10'h3]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_57 = {{_GEN_33}, {_GEN_56[{inst[14:12], inst[6:0]} == 10'h83]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_58 = {{_GEN_32}, {_GEN_57[{inst[14:12], inst[6:0]} == 10'h103]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_59 = {{_GEN_31}, {_GEN_58[{inst[14:12], inst[6:0]} == 10'h203]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_60 = {{_GEN_30}, {_GEN_59[{inst[14:12], inst[6:0]} == 10'h283]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_61 = {{_GEN_29}, {_GEN_60[{inst[14:12], inst[6:0]} == 10'h23]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_62 = {{_GEN_28}, {_GEN_61[{inst[14:12], inst[6:0]} == 10'hA3]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_63 = {{_GEN_27}, {_GEN_62[{inst[14:12], inst[6:0]} == 10'h123]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_64 = {{_GEN_26}, {_GEN_63[{inst[14:12], inst[6:0]} == 10'h13]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_65 = {{_GEN_25}, {_GEN_64[{inst[14:12], inst[6:0]} == 10'h113]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_66 = {{_GEN_24}, {_GEN_65[{inst[14:12], inst[6:0]} == 10'h193]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_67 = {{_GEN_23}, {_GEN_66[{inst[14:12], inst[6:0]} == 10'h213]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_68 = {{_GEN_22}, {_GEN_67[{inst[14:12], inst[6:0]} == 10'h313]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_69 = {{_GEN_21}, {_GEN_68[{inst[14:12], inst[6:0]} == 10'h393]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_70 = {{_GEN_20}, {_GEN_69[{inst[31:25], inst[14:12], inst[6:0]} == 17'h93]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_71 = {{_GEN_19}, {_GEN_70[{inst[31:25], inst[14:12], inst[6:0]} == 17'h293]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_72 = {{_GEN_18}, {_GEN_71[{inst[31:25], inst[14:12], inst[6:0]} == 17'h8293]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_73 = {{_GEN_17}, {_GEN_72[{inst[31:25], inst[14:12], inst[6:0]} == 17'h33]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_74 = {{_GEN_16}, {_GEN_73[{inst[31:25], inst[14:12], inst[6:0]} == 17'h8033]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_75 = {{_GEN_15}, {_GEN_74[{inst[31:25], inst[14:12], inst[6:0]} == 17'hB3]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_76 = {{_GEN_14}, {_GEN_75[{inst[31:25], inst[14:12], inst[6:0]} == 17'h133]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_77 = {{_GEN_13}, {_GEN_76[{inst[31:25], inst[14:12], inst[6:0]} == 17'h1B3]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_78 = {{_GEN_12}, {_GEN_77[{inst[31:25], inst[14:12], inst[6:0]} == 17'h233]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_79 = {{_GEN_11}, {_GEN_78[{inst[31:25], inst[14:12], inst[6:0]} == 17'h2B3]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_80 = {{_GEN_10}, {_GEN_79[{inst[31:25], inst[14:12], inst[6:0]} == 17'h82B3]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_81 = {{_GEN_9}, {_GEN_80[{inst[31:25], inst[14:12], inst[6:0]} == 17'h333]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_82 = {{_GEN}, {_GEN_81[{inst[31:25], inst[14:12], inst[6:0]} == 17'h3B3]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_83 = {{_GEN_8}, {_GEN_82[{inst[31:28], inst[19:0]} == 24'hF]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_84 = {{_GEN_7}, {_GEN_83[inst == 32'h100F]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_85 = {{_GEN_6}, {_GEN_84[{inst[14:12], inst[6:0]} == 10'hF3]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_86 = {{_GEN_5}, {_GEN_85[{inst[14:12], inst[6:0]} == 10'h173]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_87 = {{_GEN_4}, {_GEN_86[{inst[14:12], inst[6:0]} == 10'h1F3]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_88 = {{_GEN_3}, {_GEN_87[{inst[14:12], inst[6:0]} == 10'h2F3]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_89 = {{_GEN_2}, {_GEN_88[{inst[14:12], inst[6:0]} == 10'h373]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_90 = {{_GEN_1}, {_GEN_89[{inst[14:12], inst[6:0]} == 10'h3F3]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_91 = {{_GEN_1}, {_GEN_90[inst == 32'h73]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_92 = {{_GEN_0}, {_GEN_91[inst == 32'h100073]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }[1:0]
    _GEN_93 = {{_GEN}, {_GEN_92[inst == 32'h10000073]}};
  wire
    struct packed {logic [1:0] _0; logic _1; logic _2; logic [2:0] _3; logic [3:0] _4; logic [2:0] _5; logic _6; logic [1:0] _7; logic [2:0] _8; logic [1:0] _9; logic _10; logic [2:0] _11; logic _12; }
    _GEN_94 = _GEN_93[inst == 32'h10200073];
  assign pc_sel = _GEN_94._0;
  assign inst_kill = _GEN_94._6;
  assign A_sel = _GEN_94._1;
  assign B_sel = _GEN_94._2;
  assign imm_sel = _GEN_94._3;
  assign alu_op = _GEN_94._4;
  assign br_type = _GEN_94._5;
  assign st_type = _GEN_94._7;
  assign ld_type = _GEN_94._8;
  assign wb_sel = _GEN_94._9;
  assign wb_en = _GEN_94._10;
  assign csr_cmd = _GEN_94._11;
  assign illegal = _GEN_94._12;
endmodule

module Core(
  input  struct packed {logic valid; logic [31:0] data; }                                                             host_fromhost,
  input  struct packed {logic valid; struct packed {logic [31:0] data; } data; }                                      icache_resp,
                                                                                                                      dcache_resp,
  input                                                                                                               CLK,
                                                                                                                      RESET,
  output [31:0]                                                                                                       host_tohost,
  output                                                                                                              icache_abort,
  output struct packed {logic valid; struct packed {logic [31:0] addr; logic [31:0] data; logic [3:0] mask; } data; } icache_req,
  output                                                                                                              dcache_abort,
  output struct packed {logic valid; struct packed {logic [31:0] addr; logic [31:0] data; logic [3:0] mask; } data; } dcache_req
);

  wire [31:0] _Datapath_inst0_ctrl_inst;
  wire [1:0]  _Control_inst0_pc_sel;
  wire        _Control_inst0_inst_kill;
  wire        _Control_inst0_A_sel;
  wire        _Control_inst0_B_sel;
  wire [2:0]  _Control_inst0_imm_sel;
  wire [3:0]  _Control_inst0_alu_op;
  wire [2:0]  _Control_inst0_br_type;
  wire [1:0]  _Control_inst0_st_type;
  wire [2:0]  _Control_inst0_ld_type;
  wire [1:0]  _Control_inst0_wb_sel;
  wire        _Control_inst0_wb_en;
  wire [2:0]  _Control_inst0_csr_cmd;
  wire        _Control_inst0_illegal;
  Control Control_inst0 (
    .inst      (_Datapath_inst0_ctrl_inst),
    .pc_sel    (_Control_inst0_pc_sel),
    .inst_kill (_Control_inst0_inst_kill),
    .A_sel     (_Control_inst0_A_sel),
    .B_sel     (_Control_inst0_B_sel),
    .imm_sel   (_Control_inst0_imm_sel),
    .alu_op    (_Control_inst0_alu_op),
    .br_type   (_Control_inst0_br_type),
    .st_type   (_Control_inst0_st_type),
    .ld_type   (_Control_inst0_ld_type),
    .wb_sel    (_Control_inst0_wb_sel),
    .wb_en     (_Control_inst0_wb_en),
    .csr_cmd   (_Control_inst0_csr_cmd),
    .illegal   (_Control_inst0_illegal)
  );
  Datapath Datapath_inst0 (
    .host_fromhost  (host_fromhost),
    .icache_resp    (icache_resp),
    .dcache_resp    (dcache_resp),
    .ctrl_pc_sel    (_Control_inst0_pc_sel),
    .ctrl_inst_kill (_Control_inst0_inst_kill),
    .ctrl_A_sel     (_Control_inst0_A_sel),
    .ctrl_B_sel     (_Control_inst0_B_sel),
    .ctrl_imm_sel   (_Control_inst0_imm_sel),
    .ctrl_alu_op    (_Control_inst0_alu_op),
    .ctrl_br_type   (_Control_inst0_br_type),
    .ctrl_st_type   (_Control_inst0_st_type),
    .ctrl_ld_type   (_Control_inst0_ld_type),
    .ctrl_wb_sel    (_Control_inst0_wb_sel),
    .ctrl_wb_en     (_Control_inst0_wb_en),
    .ctrl_csr_cmd   (_Control_inst0_csr_cmd),
    .ctrl_illegal   (_Control_inst0_illegal),
    .CLK            (CLK),
    .RESET          (RESET),
    .host_tohost    (host_tohost),
    .icache_abort   (icache_abort),
    .icache_req     (icache_req),
    .dcache_abort   (dcache_abort),
    .dcache_req     (dcache_req),
    .ctrl_inst      (_Datapath_inst0_ctrl_inst)
  );
endmodule

module Memory(
  input  [7:0]                              RADDR,
  input                                     CLK,
                                            RE,
  input  [7:0]                              WADDR,
  input  struct packed {logic [19:0] tag; } WDATA,
  input                                     WE,
  output struct packed {logic [19:0] tag; } RDATA
);

  reg  [255:0][19:0] coreir_mem256x20_inst0;
  reg  [19:0]        read_reg;
  always_ff @(posedge CLK) begin
    if (WE)
      coreir_mem256x20_inst0[WADDR] <= WDATA.tag;
    if (RE)
      read_reg <= coreir_mem256x20_inst0[RADDR];
  end // always_ff @(posedge)
  wire struct packed {logic [19:0] tag; } _GEN;
  assign _GEN.tag = read_reg;
  assign RDATA = _GEN;
endmodule

module Memory_unq1(
  input  [7:0] RADDR,
  input        CLK,
               RE,
  input  [7:0] WADDR,
               WDATA,
  input        WE,
  output [7:0] RDATA
);

  reg [255:0][7:0] coreir_mem256x8_inst0;
  reg [7:0]        read_reg;
  always_ff @(posedge CLK) begin
    if (WE)
      coreir_mem256x8_inst0[WADDR] <= WDATA;
    if (RE)
      read_reg <= coreir_mem256x8_inst0[RADDR];
  end // always_ff @(posedge)
  assign RDATA = read_reg;
endmodule

module ArrayMaskMem(
  input  [7:0]      RADDR,
  input             CLK,
                    RE,
  input  [7:0]      WADDR,
  input  [3:0][7:0] WDATA,
  input  [3:0]      WMASK,
  input             WE,
  output [3:0][7:0] RDATA
);

  wire [7:0] _Memory_inst3_RDATA;
  wire [7:0] _Memory_inst2_RDATA;
  wire [7:0] _Memory_inst1_RDATA;
  wire [7:0] _Memory_inst0_RDATA;
  Memory_unq1 Memory_inst0 (
    .RADDR (RADDR),
    .CLK   (CLK),
    .RE    (RE),
    .WADDR (WADDR),
    .WDATA (WDATA[2'h0]),
    .WE    (WE & WMASK[0]),
    .RDATA (_Memory_inst0_RDATA)
  );
  Memory_unq1 Memory_inst1 (
    .RADDR (RADDR),
    .CLK   (CLK),
    .RE    (RE),
    .WADDR (WADDR),
    .WDATA (WDATA[2'h1]),
    .WE    (WE & WMASK[1]),
    .RDATA (_Memory_inst1_RDATA)
  );
  Memory_unq1 Memory_inst2 (
    .RADDR (RADDR),
    .CLK   (CLK),
    .RE    (RE),
    .WADDR (WADDR),
    .WDATA (WDATA[2'h2]),
    .WE    (WE & WMASK[2]),
    .RDATA (_Memory_inst2_RDATA)
  );
  Memory_unq1 Memory_inst3 (
    .RADDR (RADDR),
    .CLK   (CLK),
    .RE    (RE),
    .WADDR (WADDR),
    .WDATA (WDATA[2'h3]),
    .WE    (WE & WMASK[3]),
    .RDATA (_Memory_inst3_RDATA)
  );
  assign RDATA =
    {{_Memory_inst3_RDATA},
     {_Memory_inst2_RDATA},
     {_Memory_inst1_RDATA},
     {_Memory_inst0_RDATA}};
endmodule

module Counter(
  input  CLK,
         CE,
         RESET,
  output O,
         COUT
);

  reg Register_inst0;
  always_ff @(posedge CLK) begin
    if (RESET)
      Register_inst0 <= 1'h0;
    else begin
      if (CE)
        Register_inst0 <= Register_inst0 - 1'h1;
    end
  end // always_ff @(posedge)
  initial
    Register_inst0 = 1'h0;
  assign O = Register_inst0;
  assign COUT = Register_inst0 & CE;
endmodule

module Cache(
  input                                                                                                                                                                                                                 cpu_abort,
  input  struct packed {logic valid; struct packed {logic [31:0] addr; logic [31:0] data; logic [3:0] mask; } data; }                                                                                                   cpu_req,
  input                                                                                                                                                                                                                 nasti_aw_ready,
                                                                                                                                                                                                                        nasti_w_ready,
                                                                                                                                                                                                                        nasti_b_valid,
  input  struct packed {logic [1:0] resp; logic [4:0] id; logic user; }                                                                                                                                                 nasti_b_data,
  input                                                                                                                                                                                                                 nasti_ar_ready,
                                                                                                                                                                                                                        nasti_r_valid,
  input  struct packed {logic [1:0] resp; logic [4:0] id; logic user; logic [63:0] data; logic last; }                                                                                                                  nasti_r_data,
  input                                                                                                                                                                                                                 CLK,
                                                                                                                                                                                                                        RESET,
  output struct packed {logic valid; struct packed {logic [31:0] data; } data; }                                                                                                                                        cpu_resp,
  output                                                                                                                                                                                                                nasti_aw_valid,
  output struct packed {logic [4:0] id; logic user; logic [31:0] addr; logic [7:0] length; logic [2:0] size; logic [1:0] burst; logic lock; logic [3:0] cache; logic [2:0] prot; logic [3:0] qos; logic [3:0] region; } nasti_aw_data,
  output                                                                                                                                                                                                                nasti_w_valid,
  output struct packed {logic [4:0] id; logic [7:0] strb; logic user; logic [63:0] data; logic last; }                                                                                                                  nasti_w_data,
  output                                                                                                                                                                                                                nasti_b_ready,
                                                                                                                                                                                                                        nasti_ar_valid,
  output struct packed {logic [4:0] id; logic user; logic [31:0] addr; logic [7:0] length; logic [2:0] size; logic [1:0] burst; logic lock; logic [3:0] cache; logic [2:0] prot; logic [3:0] qos; logic [3:0] region; } nasti_ar_data,
  output                                                                                                                                                                                                                nasti_r_ready
);

  reg  [1:0][63:0]  Register_inst6;
  wire              _GEN;
  reg  [2:0]        Register_inst0;
  reg               _GEN_0;
  reg               _GEN_1;
  reg               _GEN_2;
  reg               _GEN_3;
  wire              hit;
  wire [3:0][7:0]   _ArrayMaskMem_inst3_RDATA;
  wire [3:0][7:0]   _ArrayMaskMem_inst2_RDATA;
  wire [3:0][7:0]   _ArrayMaskMem_inst1_RDATA;
  wire [3:0][7:0]   _ArrayMaskMem_inst0_RDATA;
  wire              _Counter_inst1_O;
  wire              _Counter_inst1_COUT;
  wire struct packed {logic [19:0] tag; } _Memory_inst0_RDATA;
  wire              _Counter_inst0_O;
  wire              _Counter_inst0_COUT;
  reg  [31:0]       Register_inst3;
  wire              _GEN_4 = Register_inst0 == 3'h6;
  wire              _GEN_5 = Register_inst0 == 3'h6 & _Counter_inst0_COUT;
  reg               Register_inst7;
  wire              _GEN_6 =
    Register_inst0 == 3'h2 & (hit | Register_inst7) & ~cpu_abort | _GEN_5;
  reg  [255:0]      Register_inst1;
  wire [255:0]      _GEN_7 = Register_inst1 >> Register_inst3[11:4];
  wire              _GEN_8 = Register_inst0 == 3'h1;
  wire              _GEN_9 = ~_GEN_6 & (_GEN | _GEN_8) & cpu_req.valid;
  wire struct packed {logic [19:0] tag; } _GEN_10;
  assign _GEN_10.tag = Register_inst3[31:12];
  wire struct packed {logic [19:0] tag; } wmeta = _GEN_10;
  assign hit = _GEN_7[0] & _Memory_inst0_RDATA.tag == Register_inst3[31:12];
  reg  [255:0]      Register_inst2;
  wire              aw_valid = _GEN_3;
  wire              ar_valid = _GEN_2;
  wire              b_ready = _GEN_0;
  reg  [3:0]        Register_inst5;
  reg  [2:0]        _GEN_11;
  wire [255:0]      _GEN_12 = Register_inst2 >> Register_inst3[11:4];
  wire [255:0]      _GEN_13 = Register_inst1 >> Register_inst3[11:4];
  wire              _GEN_14 = _GEN_13[0] & _GEN_12[0];
  always_comb begin
    _GEN_11 = Register_inst0;
    _GEN_3 = 1'h0;
    _GEN_2 = 1'h0;
    _GEN_1 = 1'h0;
    _GEN_0 = 1'h0;
    if (Register_inst0 == 3'h0) begin
      if (cpu_req.valid) begin
        if (|cpu_req.data.mask)
          _GEN_11 = 3'h2;
        else
          _GEN_11 = 3'h1;
      end
    end
    else if (Register_inst0 == 3'h1) begin
      if (hit) begin
        if (cpu_req.valid) begin
          if (|cpu_req.data.mask)
            _GEN_11 = 3'h2;
          else
            _GEN_11 = 3'h1;
        end
        else
          _GEN_11 = 3'h0;
      end
      else begin
        _GEN_3 = _GEN_14;
        _GEN_2 = ~_GEN_14;
        if (nasti_aw_ready & aw_valid)
          _GEN_11 = 3'h3;
        else if (nasti_ar_ready & ar_valid)
          _GEN_11 = 3'h6;
      end
    end
    else if (Register_inst0 == 3'h2) begin
      if (hit | Register_inst7 | cpu_abort)
        _GEN_11 = 3'h0;
      else begin
        _GEN_3 = _GEN_14;
        _GEN_2 = ~_GEN_14;
        if (nasti_aw_ready & aw_valid)
          _GEN_11 = 3'h3;
        else if (nasti_ar_ready & ar_valid)
          _GEN_11 = 3'h6;
      end
    end
    else if (Register_inst0 == 3'h3) begin
      _GEN_1 = 1'h1;
      if (_Counter_inst1_COUT)
        _GEN_11 = 3'h4;
    end
    else if (Register_inst0 == 3'h4) begin
      _GEN_0 = 1'h1;
      if (b_ready & nasti_b_valid)
        _GEN_11 = 3'h5;
    end
    else if (Register_inst0 == 3'h5) begin
      _GEN_2 = 1'h1;
      if (nasti_ar_ready & ar_valid)
        _GEN_11 = 3'h6;
    end
    else if (Register_inst0 == 3'h6) begin
      if (_Counter_inst0_COUT) begin
        if (|Register_inst5)
          _GEN_11 = 3'h2;
        else
          _GEN_11 = 3'h0;
      end
    end
  end // always_comb
  always_ff @(posedge CLK) begin
    if (RESET)
      Register_inst0 <= 3'h0;
    else
      Register_inst0 <= _GEN_11;
  end // always_ff @(posedge)
  assign _GEN = Register_inst0 == 3'h0;
  wire              _GEN_15 =
    _GEN | _GEN_8 & hit | Register_inst7 & Register_inst5 == 4'h0;
  reg  [31:0]       Register_inst4;
  wire [1:0][127:0] _GEN_16 =
    {{{4{Register_inst4}}}, {{nasti_r_data.data, Register_inst6[1'h0]}}};
  wire [127:0]      _GEN_17 = _GEN_16[~_GEN_5];
  wire [1:0][31:0]  _GEN_18 =
    {{{28'h0, Register_inst5} << {28'h0, Register_inst3[3:2], 2'h0}}, {32'hFFFFFFFF}};
  wire [31:0]       _GEN_19 = _GEN_18[~_GEN_5];
  reg               Register_inst8;
  reg  [15:0][7:0]  Register_inst9;
  wire [1:0]        _GEN_20 = {{1'h1}, {Register_inst1[255]}};
  wire [1:0]        _GEN_21 = {{1'h1}, {Register_inst1[254]}};
  wire [1:0]        _GEN_22 = {{1'h1}, {Register_inst1[253]}};
  wire [1:0]        _GEN_23 = {{1'h1}, {Register_inst1[252]}};
  wire [1:0]        _GEN_24 = {{1'h1}, {Register_inst1[251]}};
  wire [1:0]        _GEN_25 = {{1'h1}, {Register_inst1[250]}};
  wire [1:0]        _GEN_26 = {{1'h1}, {Register_inst1[249]}};
  wire [1:0]        _GEN_27 = {{1'h1}, {Register_inst1[248]}};
  wire [1:0]        _GEN_28 = {{1'h1}, {Register_inst1[247]}};
  wire [1:0]        _GEN_29 = {{1'h1}, {Register_inst1[246]}};
  wire [1:0]        _GEN_30 = {{1'h1}, {Register_inst1[245]}};
  wire [1:0]        _GEN_31 = {{1'h1}, {Register_inst1[244]}};
  wire [1:0]        _GEN_32 = {{1'h1}, {Register_inst1[243]}};
  wire [1:0]        _GEN_33 = {{1'h1}, {Register_inst1[242]}};
  wire [1:0]        _GEN_34 = {{1'h1}, {Register_inst1[241]}};
  wire [1:0]        _GEN_35 = {{1'h1}, {Register_inst1[240]}};
  wire [1:0]        _GEN_36 = {{1'h1}, {Register_inst1[239]}};
  wire [1:0]        _GEN_37 = {{1'h1}, {Register_inst1[238]}};
  wire [1:0]        _GEN_38 = {{1'h1}, {Register_inst1[237]}};
  wire [1:0]        _GEN_39 = {{1'h1}, {Register_inst1[236]}};
  wire [1:0]        _GEN_40 = {{1'h1}, {Register_inst1[235]}};
  wire [1:0]        _GEN_41 = {{1'h1}, {Register_inst1[234]}};
  wire [1:0]        _GEN_42 = {{1'h1}, {Register_inst1[233]}};
  wire [1:0]        _GEN_43 = {{1'h1}, {Register_inst1[232]}};
  wire [1:0]        _GEN_44 = {{1'h1}, {Register_inst1[231]}};
  wire [1:0]        _GEN_45 = {{1'h1}, {Register_inst1[230]}};
  wire [1:0]        _GEN_46 = {{1'h1}, {Register_inst1[229]}};
  wire [1:0]        _GEN_47 = {{1'h1}, {Register_inst1[228]}};
  wire [1:0]        _GEN_48 = {{1'h1}, {Register_inst1[227]}};
  wire [1:0]        _GEN_49 = {{1'h1}, {Register_inst1[226]}};
  wire [1:0]        _GEN_50 = {{1'h1}, {Register_inst1[225]}};
  wire [1:0]        _GEN_51 = {{1'h1}, {Register_inst1[224]}};
  wire [1:0]        _GEN_52 = {{1'h1}, {Register_inst1[223]}};
  wire [1:0]        _GEN_53 = {{1'h1}, {Register_inst1[222]}};
  wire [1:0]        _GEN_54 = {{1'h1}, {Register_inst1[221]}};
  wire [1:0]        _GEN_55 = {{1'h1}, {Register_inst1[220]}};
  wire [1:0]        _GEN_56 = {{1'h1}, {Register_inst1[219]}};
  wire [1:0]        _GEN_57 = {{1'h1}, {Register_inst1[218]}};
  wire [1:0]        _GEN_58 = {{1'h1}, {Register_inst1[217]}};
  wire [1:0]        _GEN_59 = {{1'h1}, {Register_inst1[216]}};
  wire [1:0]        _GEN_60 = {{1'h1}, {Register_inst1[215]}};
  wire [1:0]        _GEN_61 = {{1'h1}, {Register_inst1[214]}};
  wire [1:0]        _GEN_62 = {{1'h1}, {Register_inst1[213]}};
  wire [1:0]        _GEN_63 = {{1'h1}, {Register_inst1[212]}};
  wire [1:0]        _GEN_64 = {{1'h1}, {Register_inst1[211]}};
  wire [1:0]        _GEN_65 = {{1'h1}, {Register_inst1[210]}};
  wire [1:0]        _GEN_66 = {{1'h1}, {Register_inst1[209]}};
  wire [1:0]        _GEN_67 = {{1'h1}, {Register_inst1[208]}};
  wire [1:0]        _GEN_68 = {{1'h1}, {Register_inst1[207]}};
  wire [1:0]        _GEN_69 = {{1'h1}, {Register_inst1[206]}};
  wire [1:0]        _GEN_70 = {{1'h1}, {Register_inst1[205]}};
  wire [1:0]        _GEN_71 = {{1'h1}, {Register_inst1[204]}};
  wire [1:0]        _GEN_72 = {{1'h1}, {Register_inst1[203]}};
  wire [1:0]        _GEN_73 = {{1'h1}, {Register_inst1[202]}};
  wire [1:0]        _GEN_74 = {{1'h1}, {Register_inst1[201]}};
  wire [1:0]        _GEN_75 = {{1'h1}, {Register_inst1[200]}};
  wire [1:0]        _GEN_76 = {{1'h1}, {Register_inst1[199]}};
  wire [1:0]        _GEN_77 = {{1'h1}, {Register_inst1[198]}};
  wire [1:0]        _GEN_78 = {{1'h1}, {Register_inst1[197]}};
  wire [1:0]        _GEN_79 = {{1'h1}, {Register_inst1[196]}};
  wire [1:0]        _GEN_80 = {{1'h1}, {Register_inst1[195]}};
  wire [1:0]        _GEN_81 = {{1'h1}, {Register_inst1[194]}};
  wire [1:0]        _GEN_82 = {{1'h1}, {Register_inst1[193]}};
  wire [1:0]        _GEN_83 = {{1'h1}, {Register_inst1[192]}};
  wire [1:0]        _GEN_84 = {{1'h1}, {Register_inst1[191]}};
  wire [1:0]        _GEN_85 = {{1'h1}, {Register_inst1[190]}};
  wire [1:0]        _GEN_86 = {{1'h1}, {Register_inst1[189]}};
  wire [1:0]        _GEN_87 = {{1'h1}, {Register_inst1[188]}};
  wire [1:0]        _GEN_88 = {{1'h1}, {Register_inst1[187]}};
  wire [1:0]        _GEN_89 = {{1'h1}, {Register_inst1[186]}};
  wire [1:0]        _GEN_90 = {{1'h1}, {Register_inst1[185]}};
  wire [1:0]        _GEN_91 = {{1'h1}, {Register_inst1[184]}};
  wire [1:0]        _GEN_92 = {{1'h1}, {Register_inst1[183]}};
  wire [1:0]        _GEN_93 = {{1'h1}, {Register_inst1[182]}};
  wire [1:0]        _GEN_94 = {{1'h1}, {Register_inst1[181]}};
  wire [1:0]        _GEN_95 = {{1'h1}, {Register_inst1[180]}};
  wire [1:0]        _GEN_96 = {{1'h1}, {Register_inst1[179]}};
  wire [1:0]        _GEN_97 = {{1'h1}, {Register_inst1[178]}};
  wire [1:0]        _GEN_98 = {{1'h1}, {Register_inst1[177]}};
  wire [1:0]        _GEN_99 = {{1'h1}, {Register_inst1[176]}};
  wire [1:0]        _GEN_100 = {{1'h1}, {Register_inst1[175]}};
  wire [1:0]        _GEN_101 = {{1'h1}, {Register_inst1[174]}};
  wire [1:0]        _GEN_102 = {{1'h1}, {Register_inst1[173]}};
  wire [1:0]        _GEN_103 = {{1'h1}, {Register_inst1[172]}};
  wire [1:0]        _GEN_104 = {{1'h1}, {Register_inst1[171]}};
  wire [1:0]        _GEN_105 = {{1'h1}, {Register_inst1[170]}};
  wire [1:0]        _GEN_106 = {{1'h1}, {Register_inst1[169]}};
  wire [1:0]        _GEN_107 = {{1'h1}, {Register_inst1[168]}};
  wire [1:0]        _GEN_108 = {{1'h1}, {Register_inst1[167]}};
  wire [1:0]        _GEN_109 = {{1'h1}, {Register_inst1[166]}};
  wire [1:0]        _GEN_110 = {{1'h1}, {Register_inst1[165]}};
  wire [1:0]        _GEN_111 = {{1'h1}, {Register_inst1[164]}};
  wire [1:0]        _GEN_112 = {{1'h1}, {Register_inst1[163]}};
  wire [1:0]        _GEN_113 = {{1'h1}, {Register_inst1[162]}};
  wire [1:0]        _GEN_114 = {{1'h1}, {Register_inst1[161]}};
  wire [1:0]        _GEN_115 = {{1'h1}, {Register_inst1[160]}};
  wire [1:0]        _GEN_116 = {{1'h1}, {Register_inst1[159]}};
  wire [1:0]        _GEN_117 = {{1'h1}, {Register_inst1[158]}};
  wire [1:0]        _GEN_118 = {{1'h1}, {Register_inst1[157]}};
  wire [1:0]        _GEN_119 = {{1'h1}, {Register_inst1[156]}};
  wire [1:0]        _GEN_120 = {{1'h1}, {Register_inst1[155]}};
  wire [1:0]        _GEN_121 = {{1'h1}, {Register_inst1[154]}};
  wire [1:0]        _GEN_122 = {{1'h1}, {Register_inst1[153]}};
  wire [1:0]        _GEN_123 = {{1'h1}, {Register_inst1[152]}};
  wire [1:0]        _GEN_124 = {{1'h1}, {Register_inst1[151]}};
  wire [1:0]        _GEN_125 = {{1'h1}, {Register_inst1[150]}};
  wire [1:0]        _GEN_126 = {{1'h1}, {Register_inst1[149]}};
  wire [1:0]        _GEN_127 = {{1'h1}, {Register_inst1[148]}};
  wire [1:0]        _GEN_128 = {{1'h1}, {Register_inst1[147]}};
  wire [1:0]        _GEN_129 = {{1'h1}, {Register_inst1[146]}};
  wire [1:0]        _GEN_130 = {{1'h1}, {Register_inst1[145]}};
  wire [1:0]        _GEN_131 = {{1'h1}, {Register_inst1[144]}};
  wire [1:0]        _GEN_132 = {{1'h1}, {Register_inst1[143]}};
  wire [1:0]        _GEN_133 = {{1'h1}, {Register_inst1[142]}};
  wire [1:0]        _GEN_134 = {{1'h1}, {Register_inst1[141]}};
  wire [1:0]        _GEN_135 = {{1'h1}, {Register_inst1[140]}};
  wire [1:0]        _GEN_136 = {{1'h1}, {Register_inst1[139]}};
  wire [1:0]        _GEN_137 = {{1'h1}, {Register_inst1[138]}};
  wire [1:0]        _GEN_138 = {{1'h1}, {Register_inst1[137]}};
  wire [1:0]        _GEN_139 = {{1'h1}, {Register_inst1[136]}};
  wire [1:0]        _GEN_140 = {{1'h1}, {Register_inst1[135]}};
  wire [1:0]        _GEN_141 = {{1'h1}, {Register_inst1[134]}};
  wire [1:0]        _GEN_142 = {{1'h1}, {Register_inst1[133]}};
  wire [1:0]        _GEN_143 = {{1'h1}, {Register_inst1[132]}};
  wire [1:0]        _GEN_144 = {{1'h1}, {Register_inst1[131]}};
  wire [1:0]        _GEN_145 = {{1'h1}, {Register_inst1[130]}};
  wire [1:0]        _GEN_146 = {{1'h1}, {Register_inst1[129]}};
  wire [1:0]        _GEN_147 = {{1'h1}, {Register_inst1[128]}};
  wire [1:0]        _GEN_148 = {{1'h1}, {Register_inst1[127]}};
  wire [1:0]        _GEN_149 = {{1'h1}, {Register_inst1[126]}};
  wire [1:0]        _GEN_150 = {{1'h1}, {Register_inst1[125]}};
  wire [1:0]        _GEN_151 = {{1'h1}, {Register_inst1[124]}};
  wire [1:0]        _GEN_152 = {{1'h1}, {Register_inst1[123]}};
  wire [1:0]        _GEN_153 = {{1'h1}, {Register_inst1[122]}};
  wire [1:0]        _GEN_154 = {{1'h1}, {Register_inst1[121]}};
  wire [1:0]        _GEN_155 = {{1'h1}, {Register_inst1[120]}};
  wire [1:0]        _GEN_156 = {{1'h1}, {Register_inst1[119]}};
  wire [1:0]        _GEN_157 = {{1'h1}, {Register_inst1[118]}};
  wire [1:0]        _GEN_158 = {{1'h1}, {Register_inst1[117]}};
  wire [1:0]        _GEN_159 = {{1'h1}, {Register_inst1[116]}};
  wire [1:0]        _GEN_160 = {{1'h1}, {Register_inst1[115]}};
  wire [1:0]        _GEN_161 = {{1'h1}, {Register_inst1[114]}};
  wire [1:0]        _GEN_162 = {{1'h1}, {Register_inst1[113]}};
  wire [1:0]        _GEN_163 = {{1'h1}, {Register_inst1[112]}};
  wire [1:0]        _GEN_164 = {{1'h1}, {Register_inst1[111]}};
  wire [1:0]        _GEN_165 = {{1'h1}, {Register_inst1[110]}};
  wire [1:0]        _GEN_166 = {{1'h1}, {Register_inst1[109]}};
  wire [1:0]        _GEN_167 = {{1'h1}, {Register_inst1[108]}};
  wire [1:0]        _GEN_168 = {{1'h1}, {Register_inst1[107]}};
  wire [1:0]        _GEN_169 = {{1'h1}, {Register_inst1[106]}};
  wire [1:0]        _GEN_170 = {{1'h1}, {Register_inst1[105]}};
  wire [1:0]        _GEN_171 = {{1'h1}, {Register_inst1[104]}};
  wire [1:0]        _GEN_172 = {{1'h1}, {Register_inst1[103]}};
  wire [1:0]        _GEN_173 = {{1'h1}, {Register_inst1[102]}};
  wire [1:0]        _GEN_174 = {{1'h1}, {Register_inst1[101]}};
  wire [1:0]        _GEN_175 = {{1'h1}, {Register_inst1[100]}};
  wire [1:0]        _GEN_176 = {{1'h1}, {Register_inst1[99]}};
  wire [1:0]        _GEN_177 = {{1'h1}, {Register_inst1[98]}};
  wire [1:0]        _GEN_178 = {{1'h1}, {Register_inst1[97]}};
  wire [1:0]        _GEN_179 = {{1'h1}, {Register_inst1[96]}};
  wire [1:0]        _GEN_180 = {{1'h1}, {Register_inst1[95]}};
  wire [1:0]        _GEN_181 = {{1'h1}, {Register_inst1[94]}};
  wire [1:0]        _GEN_182 = {{1'h1}, {Register_inst1[93]}};
  wire [1:0]        _GEN_183 = {{1'h1}, {Register_inst1[92]}};
  wire [1:0]        _GEN_184 = {{1'h1}, {Register_inst1[91]}};
  wire [1:0]        _GEN_185 = {{1'h1}, {Register_inst1[90]}};
  wire [1:0]        _GEN_186 = {{1'h1}, {Register_inst1[89]}};
  wire [1:0]        _GEN_187 = {{1'h1}, {Register_inst1[88]}};
  wire [1:0]        _GEN_188 = {{1'h1}, {Register_inst1[87]}};
  wire [1:0]        _GEN_189 = {{1'h1}, {Register_inst1[86]}};
  wire [1:0]        _GEN_190 = {{1'h1}, {Register_inst1[85]}};
  wire [1:0]        _GEN_191 = {{1'h1}, {Register_inst1[84]}};
  wire [1:0]        _GEN_192 = {{1'h1}, {Register_inst1[83]}};
  wire [1:0]        _GEN_193 = {{1'h1}, {Register_inst1[82]}};
  wire [1:0]        _GEN_194 = {{1'h1}, {Register_inst1[81]}};
  wire [1:0]        _GEN_195 = {{1'h1}, {Register_inst1[80]}};
  wire [1:0]        _GEN_196 = {{1'h1}, {Register_inst1[79]}};
  wire [1:0]        _GEN_197 = {{1'h1}, {Register_inst1[78]}};
  wire [1:0]        _GEN_198 = {{1'h1}, {Register_inst1[77]}};
  wire [1:0]        _GEN_199 = {{1'h1}, {Register_inst1[76]}};
  wire [1:0]        _GEN_200 = {{1'h1}, {Register_inst1[75]}};
  wire [1:0]        _GEN_201 = {{1'h1}, {Register_inst1[74]}};
  wire [1:0]        _GEN_202 = {{1'h1}, {Register_inst1[73]}};
  wire [1:0]        _GEN_203 = {{1'h1}, {Register_inst1[72]}};
  wire [1:0]        _GEN_204 = {{1'h1}, {Register_inst1[71]}};
  wire [1:0]        _GEN_205 = {{1'h1}, {Register_inst1[70]}};
  wire [1:0]        _GEN_206 = {{1'h1}, {Register_inst1[69]}};
  wire [1:0]        _GEN_207 = {{1'h1}, {Register_inst1[68]}};
  wire [1:0]        _GEN_208 = {{1'h1}, {Register_inst1[67]}};
  wire [1:0]        _GEN_209 = {{1'h1}, {Register_inst1[66]}};
  wire [1:0]        _GEN_210 = {{1'h1}, {Register_inst1[65]}};
  wire [1:0]        _GEN_211 = {{1'h1}, {Register_inst1[64]}};
  wire [1:0]        _GEN_212 = {{1'h1}, {Register_inst1[63]}};
  wire [1:0]        _GEN_213 = {{1'h1}, {Register_inst1[62]}};
  wire [1:0]        _GEN_214 = {{1'h1}, {Register_inst1[61]}};
  wire [1:0]        _GEN_215 = {{1'h1}, {Register_inst1[60]}};
  wire [1:0]        _GEN_216 = {{1'h1}, {Register_inst1[59]}};
  wire [1:0]        _GEN_217 = {{1'h1}, {Register_inst1[58]}};
  wire [1:0]        _GEN_218 = {{1'h1}, {Register_inst1[57]}};
  wire [1:0]        _GEN_219 = {{1'h1}, {Register_inst1[56]}};
  wire [1:0]        _GEN_220 = {{1'h1}, {Register_inst1[55]}};
  wire [1:0]        _GEN_221 = {{1'h1}, {Register_inst1[54]}};
  wire [1:0]        _GEN_222 = {{1'h1}, {Register_inst1[53]}};
  wire [1:0]        _GEN_223 = {{1'h1}, {Register_inst1[52]}};
  wire [1:0]        _GEN_224 = {{1'h1}, {Register_inst1[51]}};
  wire [1:0]        _GEN_225 = {{1'h1}, {Register_inst1[50]}};
  wire [1:0]        _GEN_226 = {{1'h1}, {Register_inst1[49]}};
  wire [1:0]        _GEN_227 = {{1'h1}, {Register_inst1[48]}};
  wire [1:0]        _GEN_228 = {{1'h1}, {Register_inst1[47]}};
  wire [1:0]        _GEN_229 = {{1'h1}, {Register_inst1[46]}};
  wire [1:0]        _GEN_230 = {{1'h1}, {Register_inst1[45]}};
  wire [1:0]        _GEN_231 = {{1'h1}, {Register_inst1[44]}};
  wire [1:0]        _GEN_232 = {{1'h1}, {Register_inst1[43]}};
  wire [1:0]        _GEN_233 = {{1'h1}, {Register_inst1[42]}};
  wire [1:0]        _GEN_234 = {{1'h1}, {Register_inst1[41]}};
  wire [1:0]        _GEN_235 = {{1'h1}, {Register_inst1[40]}};
  wire [1:0]        _GEN_236 = {{1'h1}, {Register_inst1[39]}};
  wire [1:0]        _GEN_237 = {{1'h1}, {Register_inst1[38]}};
  wire [1:0]        _GEN_238 = {{1'h1}, {Register_inst1[37]}};
  wire [1:0]        _GEN_239 = {{1'h1}, {Register_inst1[36]}};
  wire [1:0]        _GEN_240 = {{1'h1}, {Register_inst1[35]}};
  wire [1:0]        _GEN_241 = {{1'h1}, {Register_inst1[34]}};
  wire [1:0]        _GEN_242 = {{1'h1}, {Register_inst1[33]}};
  wire [1:0]        _GEN_243 = {{1'h1}, {Register_inst1[32]}};
  wire [1:0]        _GEN_244 = {{1'h1}, {Register_inst1[31]}};
  wire [1:0]        _GEN_245 = {{1'h1}, {Register_inst1[30]}};
  wire [1:0]        _GEN_246 = {{1'h1}, {Register_inst1[29]}};
  wire [1:0]        _GEN_247 = {{1'h1}, {Register_inst1[28]}};
  wire [1:0]        _GEN_248 = {{1'h1}, {Register_inst1[27]}};
  wire [1:0]        _GEN_249 = {{1'h1}, {Register_inst1[26]}};
  wire [1:0]        _GEN_250 = {{1'h1}, {Register_inst1[25]}};
  wire [1:0]        _GEN_251 = {{1'h1}, {Register_inst1[24]}};
  wire [1:0]        _GEN_252 = {{1'h1}, {Register_inst1[23]}};
  wire [1:0]        _GEN_253 = {{1'h1}, {Register_inst1[22]}};
  wire [1:0]        _GEN_254 = {{1'h1}, {Register_inst1[21]}};
  wire [1:0]        _GEN_255 = {{1'h1}, {Register_inst1[20]}};
  wire [1:0]        _GEN_256 = {{1'h1}, {Register_inst1[19]}};
  wire [1:0]        _GEN_257 = {{1'h1}, {Register_inst1[18]}};
  wire [1:0]        _GEN_258 = {{1'h1}, {Register_inst1[17]}};
  wire [1:0]        _GEN_259 = {{1'h1}, {Register_inst1[16]}};
  wire [1:0]        _GEN_260 = {{1'h1}, {Register_inst1[15]}};
  wire [1:0]        _GEN_261 = {{1'h1}, {Register_inst1[14]}};
  wire [1:0]        _GEN_262 = {{1'h1}, {Register_inst1[13]}};
  wire [1:0]        _GEN_263 = {{1'h1}, {Register_inst1[12]}};
  wire [1:0]        _GEN_264 = {{1'h1}, {Register_inst1[11]}};
  wire [1:0]        _GEN_265 = {{1'h1}, {Register_inst1[10]}};
  wire [1:0]        _GEN_266 = {{1'h1}, {Register_inst1[9]}};
  wire [1:0]        _GEN_267 = {{1'h1}, {Register_inst1[8]}};
  wire [1:0]        _GEN_268 = {{1'h1}, {Register_inst1[7]}};
  wire [1:0]        _GEN_269 = {{1'h1}, {Register_inst1[6]}};
  wire [1:0]        _GEN_270 = {{1'h1}, {Register_inst1[5]}};
  wire [1:0]        _GEN_271 = {{1'h1}, {Register_inst1[4]}};
  wire [1:0]        _GEN_272 = {{1'h1}, {Register_inst1[3]}};
  wire [1:0]        _GEN_273 = {{1'h1}, {Register_inst1[2]}};
  wire [1:0]        _GEN_274 = {{1'h1}, {Register_inst1[1]}};
  wire [1:0]        _GEN_275 = {{1'h1}, {Register_inst1[0]}};
  wire [255:0]      _GEN_276 =
    {_GEN_20[&(Register_inst3[11:4])],
     _GEN_21[Register_inst3[11:4] == 8'hFE],
     _GEN_22[Register_inst3[11:4] == 8'hFD],
     _GEN_23[Register_inst3[11:4] == 8'hFC],
     _GEN_24[Register_inst3[11:4] == 8'hFB],
     _GEN_25[Register_inst3[11:4] == 8'hFA],
     _GEN_26[Register_inst3[11:4] == 8'hF9],
     _GEN_27[Register_inst3[11:4] == 8'hF8],
     _GEN_28[Register_inst3[11:4] == 8'hF7],
     _GEN_29[Register_inst3[11:4] == 8'hF6],
     _GEN_30[Register_inst3[11:4] == 8'hF5],
     _GEN_31[Register_inst3[11:4] == 8'hF4],
     _GEN_32[Register_inst3[11:4] == 8'hF3],
     _GEN_33[Register_inst3[11:4] == 8'hF2],
     _GEN_34[Register_inst3[11:4] == 8'hF1],
     _GEN_35[Register_inst3[11:4] == 8'hF0],
     _GEN_36[Register_inst3[11:4] == 8'hEF],
     _GEN_37[Register_inst3[11:4] == 8'hEE],
     _GEN_38[Register_inst3[11:4] == 8'hED],
     _GEN_39[Register_inst3[11:4] == 8'hEC],
     _GEN_40[Register_inst3[11:4] == 8'hEB],
     _GEN_41[Register_inst3[11:4] == 8'hEA],
     _GEN_42[Register_inst3[11:4] == 8'hE9],
     _GEN_43[Register_inst3[11:4] == 8'hE8],
     _GEN_44[Register_inst3[11:4] == 8'hE7],
     _GEN_45[Register_inst3[11:4] == 8'hE6],
     _GEN_46[Register_inst3[11:4] == 8'hE5],
     _GEN_47[Register_inst3[11:4] == 8'hE4],
     _GEN_48[Register_inst3[11:4] == 8'hE3],
     _GEN_49[Register_inst3[11:4] == 8'hE2],
     _GEN_50[Register_inst3[11:4] == 8'hE1],
     _GEN_51[Register_inst3[11:4] == 8'hE0],
     _GEN_52[Register_inst3[11:4] == 8'hDF],
     _GEN_53[Register_inst3[11:4] == 8'hDE],
     _GEN_54[Register_inst3[11:4] == 8'hDD],
     _GEN_55[Register_inst3[11:4] == 8'hDC],
     _GEN_56[Register_inst3[11:4] == 8'hDB],
     _GEN_57[Register_inst3[11:4] == 8'hDA],
     _GEN_58[Register_inst3[11:4] == 8'hD9],
     _GEN_59[Register_inst3[11:4] == 8'hD8],
     _GEN_60[Register_inst3[11:4] == 8'hD7],
     _GEN_61[Register_inst3[11:4] == 8'hD6],
     _GEN_62[Register_inst3[11:4] == 8'hD5],
     _GEN_63[Register_inst3[11:4] == 8'hD4],
     _GEN_64[Register_inst3[11:4] == 8'hD3],
     _GEN_65[Register_inst3[11:4] == 8'hD2],
     _GEN_66[Register_inst3[11:4] == 8'hD1],
     _GEN_67[Register_inst3[11:4] == 8'hD0],
     _GEN_68[Register_inst3[11:4] == 8'hCF],
     _GEN_69[Register_inst3[11:4] == 8'hCE],
     _GEN_70[Register_inst3[11:4] == 8'hCD],
     _GEN_71[Register_inst3[11:4] == 8'hCC],
     _GEN_72[Register_inst3[11:4] == 8'hCB],
     _GEN_73[Register_inst3[11:4] == 8'hCA],
     _GEN_74[Register_inst3[11:4] == 8'hC9],
     _GEN_75[Register_inst3[11:4] == 8'hC8],
     _GEN_76[Register_inst3[11:4] == 8'hC7],
     _GEN_77[Register_inst3[11:4] == 8'hC6],
     _GEN_78[Register_inst3[11:4] == 8'hC5],
     _GEN_79[Register_inst3[11:4] == 8'hC4],
     _GEN_80[Register_inst3[11:4] == 8'hC3],
     _GEN_81[Register_inst3[11:4] == 8'hC2],
     _GEN_82[Register_inst3[11:4] == 8'hC1],
     _GEN_83[Register_inst3[11:4] == 8'hC0],
     _GEN_84[Register_inst3[11:4] == 8'hBF],
     _GEN_85[Register_inst3[11:4] == 8'hBE],
     _GEN_86[Register_inst3[11:4] == 8'hBD],
     _GEN_87[Register_inst3[11:4] == 8'hBC],
     _GEN_88[Register_inst3[11:4] == 8'hBB],
     _GEN_89[Register_inst3[11:4] == 8'hBA],
     _GEN_90[Register_inst3[11:4] == 8'hB9],
     _GEN_91[Register_inst3[11:4] == 8'hB8],
     _GEN_92[Register_inst3[11:4] == 8'hB7],
     _GEN_93[Register_inst3[11:4] == 8'hB6],
     _GEN_94[Register_inst3[11:4] == 8'hB5],
     _GEN_95[Register_inst3[11:4] == 8'hB4],
     _GEN_96[Register_inst3[11:4] == 8'hB3],
     _GEN_97[Register_inst3[11:4] == 8'hB2],
     _GEN_98[Register_inst3[11:4] == 8'hB1],
     _GEN_99[Register_inst3[11:4] == 8'hB0],
     _GEN_100[Register_inst3[11:4] == 8'hAF],
     _GEN_101[Register_inst3[11:4] == 8'hAE],
     _GEN_102[Register_inst3[11:4] == 8'hAD],
     _GEN_103[Register_inst3[11:4] == 8'hAC],
     _GEN_104[Register_inst3[11:4] == 8'hAB],
     _GEN_105[Register_inst3[11:4] == 8'hAA],
     _GEN_106[Register_inst3[11:4] == 8'hA9],
     _GEN_107[Register_inst3[11:4] == 8'hA8],
     _GEN_108[Register_inst3[11:4] == 8'hA7],
     _GEN_109[Register_inst3[11:4] == 8'hA6],
     _GEN_110[Register_inst3[11:4] == 8'hA5],
     _GEN_111[Register_inst3[11:4] == 8'hA4],
     _GEN_112[Register_inst3[11:4] == 8'hA3],
     _GEN_113[Register_inst3[11:4] == 8'hA2],
     _GEN_114[Register_inst3[11:4] == 8'hA1],
     _GEN_115[Register_inst3[11:4] == 8'hA0],
     _GEN_116[Register_inst3[11:4] == 8'h9F],
     _GEN_117[Register_inst3[11:4] == 8'h9E],
     _GEN_118[Register_inst3[11:4] == 8'h9D],
     _GEN_119[Register_inst3[11:4] == 8'h9C],
     _GEN_120[Register_inst3[11:4] == 8'h9B],
     _GEN_121[Register_inst3[11:4] == 8'h9A],
     _GEN_122[Register_inst3[11:4] == 8'h99],
     _GEN_123[Register_inst3[11:4] == 8'h98],
     _GEN_124[Register_inst3[11:4] == 8'h97],
     _GEN_125[Register_inst3[11:4] == 8'h96],
     _GEN_126[Register_inst3[11:4] == 8'h95],
     _GEN_127[Register_inst3[11:4] == 8'h94],
     _GEN_128[Register_inst3[11:4] == 8'h93],
     _GEN_129[Register_inst3[11:4] == 8'h92],
     _GEN_130[Register_inst3[11:4] == 8'h91],
     _GEN_131[Register_inst3[11:4] == 8'h90],
     _GEN_132[Register_inst3[11:4] == 8'h8F],
     _GEN_133[Register_inst3[11:4] == 8'h8E],
     _GEN_134[Register_inst3[11:4] == 8'h8D],
     _GEN_135[Register_inst3[11:4] == 8'h8C],
     _GEN_136[Register_inst3[11:4] == 8'h8B],
     _GEN_137[Register_inst3[11:4] == 8'h8A],
     _GEN_138[Register_inst3[11:4] == 8'h89],
     _GEN_139[Register_inst3[11:4] == 8'h88],
     _GEN_140[Register_inst3[11:4] == 8'h87],
     _GEN_141[Register_inst3[11:4] == 8'h86],
     _GEN_142[Register_inst3[11:4] == 8'h85],
     _GEN_143[Register_inst3[11:4] == 8'h84],
     _GEN_144[Register_inst3[11:4] == 8'h83],
     _GEN_145[Register_inst3[11:4] == 8'h82],
     _GEN_146[Register_inst3[11:4] == 8'h81],
     _GEN_147[Register_inst3[11:4] == 8'h80],
     _GEN_148[Register_inst3[11:4] == 8'h7F],
     _GEN_149[Register_inst3[11:4] == 8'h7E],
     _GEN_150[Register_inst3[11:4] == 8'h7D],
     _GEN_151[Register_inst3[11:4] == 8'h7C],
     _GEN_152[Register_inst3[11:4] == 8'h7B],
     _GEN_153[Register_inst3[11:4] == 8'h7A],
     _GEN_154[Register_inst3[11:4] == 8'h79],
     _GEN_155[Register_inst3[11:4] == 8'h78],
     _GEN_156[Register_inst3[11:4] == 8'h77],
     _GEN_157[Register_inst3[11:4] == 8'h76],
     _GEN_158[Register_inst3[11:4] == 8'h75],
     _GEN_159[Register_inst3[11:4] == 8'h74],
     _GEN_160[Register_inst3[11:4] == 8'h73],
     _GEN_161[Register_inst3[11:4] == 8'h72],
     _GEN_162[Register_inst3[11:4] == 8'h71],
     _GEN_163[Register_inst3[11:4] == 8'h70],
     _GEN_164[Register_inst3[11:4] == 8'h6F],
     _GEN_165[Register_inst3[11:4] == 8'h6E],
     _GEN_166[Register_inst3[11:4] == 8'h6D],
     _GEN_167[Register_inst3[11:4] == 8'h6C],
     _GEN_168[Register_inst3[11:4] == 8'h6B],
     _GEN_169[Register_inst3[11:4] == 8'h6A],
     _GEN_170[Register_inst3[11:4] == 8'h69],
     _GEN_171[Register_inst3[11:4] == 8'h68],
     _GEN_172[Register_inst3[11:4] == 8'h67],
     _GEN_173[Register_inst3[11:4] == 8'h66],
     _GEN_174[Register_inst3[11:4] == 8'h65],
     _GEN_175[Register_inst3[11:4] == 8'h64],
     _GEN_176[Register_inst3[11:4] == 8'h63],
     _GEN_177[Register_inst3[11:4] == 8'h62],
     _GEN_178[Register_inst3[11:4] == 8'h61],
     _GEN_179[Register_inst3[11:4] == 8'h60],
     _GEN_180[Register_inst3[11:4] == 8'h5F],
     _GEN_181[Register_inst3[11:4] == 8'h5E],
     _GEN_182[Register_inst3[11:4] == 8'h5D],
     _GEN_183[Register_inst3[11:4] == 8'h5C],
     _GEN_184[Register_inst3[11:4] == 8'h5B],
     _GEN_185[Register_inst3[11:4] == 8'h5A],
     _GEN_186[Register_inst3[11:4] == 8'h59],
     _GEN_187[Register_inst3[11:4] == 8'h58],
     _GEN_188[Register_inst3[11:4] == 8'h57],
     _GEN_189[Register_inst3[11:4] == 8'h56],
     _GEN_190[Register_inst3[11:4] == 8'h55],
     _GEN_191[Register_inst3[11:4] == 8'h54],
     _GEN_192[Register_inst3[11:4] == 8'h53],
     _GEN_193[Register_inst3[11:4] == 8'h52],
     _GEN_194[Register_inst3[11:4] == 8'h51],
     _GEN_195[Register_inst3[11:4] == 8'h50],
     _GEN_196[Register_inst3[11:4] == 8'h4F],
     _GEN_197[Register_inst3[11:4] == 8'h4E],
     _GEN_198[Register_inst3[11:4] == 8'h4D],
     _GEN_199[Register_inst3[11:4] == 8'h4C],
     _GEN_200[Register_inst3[11:4] == 8'h4B],
     _GEN_201[Register_inst3[11:4] == 8'h4A],
     _GEN_202[Register_inst3[11:4] == 8'h49],
     _GEN_203[Register_inst3[11:4] == 8'h48],
     _GEN_204[Register_inst3[11:4] == 8'h47],
     _GEN_205[Register_inst3[11:4] == 8'h46],
     _GEN_206[Register_inst3[11:4] == 8'h45],
     _GEN_207[Register_inst3[11:4] == 8'h44],
     _GEN_208[Register_inst3[11:4] == 8'h43],
     _GEN_209[Register_inst3[11:4] == 8'h42],
     _GEN_210[Register_inst3[11:4] == 8'h41],
     _GEN_211[Register_inst3[11:4] == 8'h40],
     _GEN_212[Register_inst3[11:4] == 8'h3F],
     _GEN_213[Register_inst3[11:4] == 8'h3E],
     _GEN_214[Register_inst3[11:4] == 8'h3D],
     _GEN_215[Register_inst3[11:4] == 8'h3C],
     _GEN_216[Register_inst3[11:4] == 8'h3B],
     _GEN_217[Register_inst3[11:4] == 8'h3A],
     _GEN_218[Register_inst3[11:4] == 8'h39],
     _GEN_219[Register_inst3[11:4] == 8'h38],
     _GEN_220[Register_inst3[11:4] == 8'h37],
     _GEN_221[Register_inst3[11:4] == 8'h36],
     _GEN_222[Register_inst3[11:4] == 8'h35],
     _GEN_223[Register_inst3[11:4] == 8'h34],
     _GEN_224[Register_inst3[11:4] == 8'h33],
     _GEN_225[Register_inst3[11:4] == 8'h32],
     _GEN_226[Register_inst3[11:4] == 8'h31],
     _GEN_227[Register_inst3[11:4] == 8'h30],
     _GEN_228[Register_inst3[11:4] == 8'h2F],
     _GEN_229[Register_inst3[11:4] == 8'h2E],
     _GEN_230[Register_inst3[11:4] == 8'h2D],
     _GEN_231[Register_inst3[11:4] == 8'h2C],
     _GEN_232[Register_inst3[11:4] == 8'h2B],
     _GEN_233[Register_inst3[11:4] == 8'h2A],
     _GEN_234[Register_inst3[11:4] == 8'h29],
     _GEN_235[Register_inst3[11:4] == 8'h28],
     _GEN_236[Register_inst3[11:4] == 8'h27],
     _GEN_237[Register_inst3[11:4] == 8'h26],
     _GEN_238[Register_inst3[11:4] == 8'h25],
     _GEN_239[Register_inst3[11:4] == 8'h24],
     _GEN_240[Register_inst3[11:4] == 8'h23],
     _GEN_241[Register_inst3[11:4] == 8'h22],
     _GEN_242[Register_inst3[11:4] == 8'h21],
     _GEN_243[Register_inst3[11:4] == 8'h20],
     _GEN_244[Register_inst3[11:4] == 8'h1F],
     _GEN_245[Register_inst3[11:4] == 8'h1E],
     _GEN_246[Register_inst3[11:4] == 8'h1D],
     _GEN_247[Register_inst3[11:4] == 8'h1C],
     _GEN_248[Register_inst3[11:4] == 8'h1B],
     _GEN_249[Register_inst3[11:4] == 8'h1A],
     _GEN_250[Register_inst3[11:4] == 8'h19],
     _GEN_251[Register_inst3[11:4] == 8'h18],
     _GEN_252[Register_inst3[11:4] == 8'h17],
     _GEN_253[Register_inst3[11:4] == 8'h16],
     _GEN_254[Register_inst3[11:4] == 8'h15],
     _GEN_255[Register_inst3[11:4] == 8'h14],
     _GEN_256[Register_inst3[11:4] == 8'h13],
     _GEN_257[Register_inst3[11:4] == 8'h12],
     _GEN_258[Register_inst3[11:4] == 8'h11],
     _GEN_259[Register_inst3[11:4] == 8'h10],
     _GEN_260[Register_inst3[11:4] == 8'hF],
     _GEN_261[Register_inst3[11:4] == 8'hE],
     _GEN_262[Register_inst3[11:4] == 8'hD],
     _GEN_263[Register_inst3[11:4] == 8'hC],
     _GEN_264[Register_inst3[11:4] == 8'hB],
     _GEN_265[Register_inst3[11:4] == 8'hA],
     _GEN_266[Register_inst3[11:4] == 8'h9],
     _GEN_267[Register_inst3[11:4] == 8'h8],
     _GEN_268[Register_inst3[11:4] == 8'h7],
     _GEN_269[Register_inst3[11:4] == 8'h6],
     _GEN_270[Register_inst3[11:4] == 8'h5],
     _GEN_271[Register_inst3[11:4] == 8'h4],
     _GEN_272[Register_inst3[11:4] == 8'h3],
     _GEN_273[Register_inst3[11:4] == 8'h2],
     _GEN_274[Register_inst3[11:4] == 8'h1],
     _GEN_275[Register_inst3[11:4] == 8'h0]};
  wire [1:0]        _GEN_277 = {{~_GEN_5}, {Register_inst2[255]}};
  wire [1:0]        _GEN_278 = {{~_GEN_5}, {Register_inst2[254]}};
  wire [1:0]        _GEN_279 = {{~_GEN_5}, {Register_inst2[253]}};
  wire [1:0]        _GEN_280 = {{~_GEN_5}, {Register_inst2[252]}};
  wire [1:0]        _GEN_281 = {{~_GEN_5}, {Register_inst2[251]}};
  wire [1:0]        _GEN_282 = {{~_GEN_5}, {Register_inst2[250]}};
  wire [1:0]        _GEN_283 = {{~_GEN_5}, {Register_inst2[249]}};
  wire [1:0]        _GEN_284 = {{~_GEN_5}, {Register_inst2[248]}};
  wire [1:0]        _GEN_285 = {{~_GEN_5}, {Register_inst2[247]}};
  wire [1:0]        _GEN_286 = {{~_GEN_5}, {Register_inst2[246]}};
  wire [1:0]        _GEN_287 = {{~_GEN_5}, {Register_inst2[245]}};
  wire [1:0]        _GEN_288 = {{~_GEN_5}, {Register_inst2[244]}};
  wire [1:0]        _GEN_289 = {{~_GEN_5}, {Register_inst2[243]}};
  wire [1:0]        _GEN_290 = {{~_GEN_5}, {Register_inst2[242]}};
  wire [1:0]        _GEN_291 = {{~_GEN_5}, {Register_inst2[241]}};
  wire [1:0]        _GEN_292 = {{~_GEN_5}, {Register_inst2[240]}};
  wire [1:0]        _GEN_293 = {{~_GEN_5}, {Register_inst2[239]}};
  wire [1:0]        _GEN_294 = {{~_GEN_5}, {Register_inst2[238]}};
  wire [1:0]        _GEN_295 = {{~_GEN_5}, {Register_inst2[237]}};
  wire [1:0]        _GEN_296 = {{~_GEN_5}, {Register_inst2[236]}};
  wire [1:0]        _GEN_297 = {{~_GEN_5}, {Register_inst2[235]}};
  wire [1:0]        _GEN_298 = {{~_GEN_5}, {Register_inst2[234]}};
  wire [1:0]        _GEN_299 = {{~_GEN_5}, {Register_inst2[233]}};
  wire [1:0]        _GEN_300 = {{~_GEN_5}, {Register_inst2[232]}};
  wire [1:0]        _GEN_301 = {{~_GEN_5}, {Register_inst2[231]}};
  wire [1:0]        _GEN_302 = {{~_GEN_5}, {Register_inst2[230]}};
  wire [1:0]        _GEN_303 = {{~_GEN_5}, {Register_inst2[229]}};
  wire [1:0]        _GEN_304 = {{~_GEN_5}, {Register_inst2[228]}};
  wire [1:0]        _GEN_305 = {{~_GEN_5}, {Register_inst2[227]}};
  wire [1:0]        _GEN_306 = {{~_GEN_5}, {Register_inst2[226]}};
  wire [1:0]        _GEN_307 = {{~_GEN_5}, {Register_inst2[225]}};
  wire [1:0]        _GEN_308 = {{~_GEN_5}, {Register_inst2[224]}};
  wire [1:0]        _GEN_309 = {{~_GEN_5}, {Register_inst2[223]}};
  wire [1:0]        _GEN_310 = {{~_GEN_5}, {Register_inst2[222]}};
  wire [1:0]        _GEN_311 = {{~_GEN_5}, {Register_inst2[221]}};
  wire [1:0]        _GEN_312 = {{~_GEN_5}, {Register_inst2[220]}};
  wire [1:0]        _GEN_313 = {{~_GEN_5}, {Register_inst2[219]}};
  wire [1:0]        _GEN_314 = {{~_GEN_5}, {Register_inst2[218]}};
  wire [1:0]        _GEN_315 = {{~_GEN_5}, {Register_inst2[217]}};
  wire [1:0]        _GEN_316 = {{~_GEN_5}, {Register_inst2[216]}};
  wire [1:0]        _GEN_317 = {{~_GEN_5}, {Register_inst2[215]}};
  wire [1:0]        _GEN_318 = {{~_GEN_5}, {Register_inst2[214]}};
  wire [1:0]        _GEN_319 = {{~_GEN_5}, {Register_inst2[213]}};
  wire [1:0]        _GEN_320 = {{~_GEN_5}, {Register_inst2[212]}};
  wire [1:0]        _GEN_321 = {{~_GEN_5}, {Register_inst2[211]}};
  wire [1:0]        _GEN_322 = {{~_GEN_5}, {Register_inst2[210]}};
  wire [1:0]        _GEN_323 = {{~_GEN_5}, {Register_inst2[209]}};
  wire [1:0]        _GEN_324 = {{~_GEN_5}, {Register_inst2[208]}};
  wire [1:0]        _GEN_325 = {{~_GEN_5}, {Register_inst2[207]}};
  wire [1:0]        _GEN_326 = {{~_GEN_5}, {Register_inst2[206]}};
  wire [1:0]        _GEN_327 = {{~_GEN_5}, {Register_inst2[205]}};
  wire [1:0]        _GEN_328 = {{~_GEN_5}, {Register_inst2[204]}};
  wire [1:0]        _GEN_329 = {{~_GEN_5}, {Register_inst2[203]}};
  wire [1:0]        _GEN_330 = {{~_GEN_5}, {Register_inst2[202]}};
  wire [1:0]        _GEN_331 = {{~_GEN_5}, {Register_inst2[201]}};
  wire [1:0]        _GEN_332 = {{~_GEN_5}, {Register_inst2[200]}};
  wire [1:0]        _GEN_333 = {{~_GEN_5}, {Register_inst2[199]}};
  wire [1:0]        _GEN_334 = {{~_GEN_5}, {Register_inst2[198]}};
  wire [1:0]        _GEN_335 = {{~_GEN_5}, {Register_inst2[197]}};
  wire [1:0]        _GEN_336 = {{~_GEN_5}, {Register_inst2[196]}};
  wire [1:0]        _GEN_337 = {{~_GEN_5}, {Register_inst2[195]}};
  wire [1:0]        _GEN_338 = {{~_GEN_5}, {Register_inst2[194]}};
  wire [1:0]        _GEN_339 = {{~_GEN_5}, {Register_inst2[193]}};
  wire [1:0]        _GEN_340 = {{~_GEN_5}, {Register_inst2[192]}};
  wire [1:0]        _GEN_341 = {{~_GEN_5}, {Register_inst2[191]}};
  wire [1:0]        _GEN_342 = {{~_GEN_5}, {Register_inst2[190]}};
  wire [1:0]        _GEN_343 = {{~_GEN_5}, {Register_inst2[189]}};
  wire [1:0]        _GEN_344 = {{~_GEN_5}, {Register_inst2[188]}};
  wire [1:0]        _GEN_345 = {{~_GEN_5}, {Register_inst2[187]}};
  wire [1:0]        _GEN_346 = {{~_GEN_5}, {Register_inst2[186]}};
  wire [1:0]        _GEN_347 = {{~_GEN_5}, {Register_inst2[185]}};
  wire [1:0]        _GEN_348 = {{~_GEN_5}, {Register_inst2[184]}};
  wire [1:0]        _GEN_349 = {{~_GEN_5}, {Register_inst2[183]}};
  wire [1:0]        _GEN_350 = {{~_GEN_5}, {Register_inst2[182]}};
  wire [1:0]        _GEN_351 = {{~_GEN_5}, {Register_inst2[181]}};
  wire [1:0]        _GEN_352 = {{~_GEN_5}, {Register_inst2[180]}};
  wire [1:0]        _GEN_353 = {{~_GEN_5}, {Register_inst2[179]}};
  wire [1:0]        _GEN_354 = {{~_GEN_5}, {Register_inst2[178]}};
  wire [1:0]        _GEN_355 = {{~_GEN_5}, {Register_inst2[177]}};
  wire [1:0]        _GEN_356 = {{~_GEN_5}, {Register_inst2[176]}};
  wire [1:0]        _GEN_357 = {{~_GEN_5}, {Register_inst2[175]}};
  wire [1:0]        _GEN_358 = {{~_GEN_5}, {Register_inst2[174]}};
  wire [1:0]        _GEN_359 = {{~_GEN_5}, {Register_inst2[173]}};
  wire [1:0]        _GEN_360 = {{~_GEN_5}, {Register_inst2[172]}};
  wire [1:0]        _GEN_361 = {{~_GEN_5}, {Register_inst2[171]}};
  wire [1:0]        _GEN_362 = {{~_GEN_5}, {Register_inst2[170]}};
  wire [1:0]        _GEN_363 = {{~_GEN_5}, {Register_inst2[169]}};
  wire [1:0]        _GEN_364 = {{~_GEN_5}, {Register_inst2[168]}};
  wire [1:0]        _GEN_365 = {{~_GEN_5}, {Register_inst2[167]}};
  wire [1:0]        _GEN_366 = {{~_GEN_5}, {Register_inst2[166]}};
  wire [1:0]        _GEN_367 = {{~_GEN_5}, {Register_inst2[165]}};
  wire [1:0]        _GEN_368 = {{~_GEN_5}, {Register_inst2[164]}};
  wire [1:0]        _GEN_369 = {{~_GEN_5}, {Register_inst2[163]}};
  wire [1:0]        _GEN_370 = {{~_GEN_5}, {Register_inst2[162]}};
  wire [1:0]        _GEN_371 = {{~_GEN_5}, {Register_inst2[161]}};
  wire [1:0]        _GEN_372 = {{~_GEN_5}, {Register_inst2[160]}};
  wire [1:0]        _GEN_373 = {{~_GEN_5}, {Register_inst2[159]}};
  wire [1:0]        _GEN_374 = {{~_GEN_5}, {Register_inst2[158]}};
  wire [1:0]        _GEN_375 = {{~_GEN_5}, {Register_inst2[157]}};
  wire [1:0]        _GEN_376 = {{~_GEN_5}, {Register_inst2[156]}};
  wire [1:0]        _GEN_377 = {{~_GEN_5}, {Register_inst2[155]}};
  wire [1:0]        _GEN_378 = {{~_GEN_5}, {Register_inst2[154]}};
  wire [1:0]        _GEN_379 = {{~_GEN_5}, {Register_inst2[153]}};
  wire [1:0]        _GEN_380 = {{~_GEN_5}, {Register_inst2[152]}};
  wire [1:0]        _GEN_381 = {{~_GEN_5}, {Register_inst2[151]}};
  wire [1:0]        _GEN_382 = {{~_GEN_5}, {Register_inst2[150]}};
  wire [1:0]        _GEN_383 = {{~_GEN_5}, {Register_inst2[149]}};
  wire [1:0]        _GEN_384 = {{~_GEN_5}, {Register_inst2[148]}};
  wire [1:0]        _GEN_385 = {{~_GEN_5}, {Register_inst2[147]}};
  wire [1:0]        _GEN_386 = {{~_GEN_5}, {Register_inst2[146]}};
  wire [1:0]        _GEN_387 = {{~_GEN_5}, {Register_inst2[145]}};
  wire [1:0]        _GEN_388 = {{~_GEN_5}, {Register_inst2[144]}};
  wire [1:0]        _GEN_389 = {{~_GEN_5}, {Register_inst2[143]}};
  wire [1:0]        _GEN_390 = {{~_GEN_5}, {Register_inst2[142]}};
  wire [1:0]        _GEN_391 = {{~_GEN_5}, {Register_inst2[141]}};
  wire [1:0]        _GEN_392 = {{~_GEN_5}, {Register_inst2[140]}};
  wire [1:0]        _GEN_393 = {{~_GEN_5}, {Register_inst2[139]}};
  wire [1:0]        _GEN_394 = {{~_GEN_5}, {Register_inst2[138]}};
  wire [1:0]        _GEN_395 = {{~_GEN_5}, {Register_inst2[137]}};
  wire [1:0]        _GEN_396 = {{~_GEN_5}, {Register_inst2[136]}};
  wire [1:0]        _GEN_397 = {{~_GEN_5}, {Register_inst2[135]}};
  wire [1:0]        _GEN_398 = {{~_GEN_5}, {Register_inst2[134]}};
  wire [1:0]        _GEN_399 = {{~_GEN_5}, {Register_inst2[133]}};
  wire [1:0]        _GEN_400 = {{~_GEN_5}, {Register_inst2[132]}};
  wire [1:0]        _GEN_401 = {{~_GEN_5}, {Register_inst2[131]}};
  wire [1:0]        _GEN_402 = {{~_GEN_5}, {Register_inst2[130]}};
  wire [1:0]        _GEN_403 = {{~_GEN_5}, {Register_inst2[129]}};
  wire [1:0]        _GEN_404 = {{~_GEN_5}, {Register_inst2[128]}};
  wire [1:0]        _GEN_405 = {{~_GEN_5}, {Register_inst2[127]}};
  wire [1:0]        _GEN_406 = {{~_GEN_5}, {Register_inst2[126]}};
  wire [1:0]        _GEN_407 = {{~_GEN_5}, {Register_inst2[125]}};
  wire [1:0]        _GEN_408 = {{~_GEN_5}, {Register_inst2[124]}};
  wire [1:0]        _GEN_409 = {{~_GEN_5}, {Register_inst2[123]}};
  wire [1:0]        _GEN_410 = {{~_GEN_5}, {Register_inst2[122]}};
  wire [1:0]        _GEN_411 = {{~_GEN_5}, {Register_inst2[121]}};
  wire [1:0]        _GEN_412 = {{~_GEN_5}, {Register_inst2[120]}};
  wire [1:0]        _GEN_413 = {{~_GEN_5}, {Register_inst2[119]}};
  wire [1:0]        _GEN_414 = {{~_GEN_5}, {Register_inst2[118]}};
  wire [1:0]        _GEN_415 = {{~_GEN_5}, {Register_inst2[117]}};
  wire [1:0]        _GEN_416 = {{~_GEN_5}, {Register_inst2[116]}};
  wire [1:0]        _GEN_417 = {{~_GEN_5}, {Register_inst2[115]}};
  wire [1:0]        _GEN_418 = {{~_GEN_5}, {Register_inst2[114]}};
  wire [1:0]        _GEN_419 = {{~_GEN_5}, {Register_inst2[113]}};
  wire [1:0]        _GEN_420 = {{~_GEN_5}, {Register_inst2[112]}};
  wire [1:0]        _GEN_421 = {{~_GEN_5}, {Register_inst2[111]}};
  wire [1:0]        _GEN_422 = {{~_GEN_5}, {Register_inst2[110]}};
  wire [1:0]        _GEN_423 = {{~_GEN_5}, {Register_inst2[109]}};
  wire [1:0]        _GEN_424 = {{~_GEN_5}, {Register_inst2[108]}};
  wire [1:0]        _GEN_425 = {{~_GEN_5}, {Register_inst2[107]}};
  wire [1:0]        _GEN_426 = {{~_GEN_5}, {Register_inst2[106]}};
  wire [1:0]        _GEN_427 = {{~_GEN_5}, {Register_inst2[105]}};
  wire [1:0]        _GEN_428 = {{~_GEN_5}, {Register_inst2[104]}};
  wire [1:0]        _GEN_429 = {{~_GEN_5}, {Register_inst2[103]}};
  wire [1:0]        _GEN_430 = {{~_GEN_5}, {Register_inst2[102]}};
  wire [1:0]        _GEN_431 = {{~_GEN_5}, {Register_inst2[101]}};
  wire [1:0]        _GEN_432 = {{~_GEN_5}, {Register_inst2[100]}};
  wire [1:0]        _GEN_433 = {{~_GEN_5}, {Register_inst2[99]}};
  wire [1:0]        _GEN_434 = {{~_GEN_5}, {Register_inst2[98]}};
  wire [1:0]        _GEN_435 = {{~_GEN_5}, {Register_inst2[97]}};
  wire [1:0]        _GEN_436 = {{~_GEN_5}, {Register_inst2[96]}};
  wire [1:0]        _GEN_437 = {{~_GEN_5}, {Register_inst2[95]}};
  wire [1:0]        _GEN_438 = {{~_GEN_5}, {Register_inst2[94]}};
  wire [1:0]        _GEN_439 = {{~_GEN_5}, {Register_inst2[93]}};
  wire [1:0]        _GEN_440 = {{~_GEN_5}, {Register_inst2[92]}};
  wire [1:0]        _GEN_441 = {{~_GEN_5}, {Register_inst2[91]}};
  wire [1:0]        _GEN_442 = {{~_GEN_5}, {Register_inst2[90]}};
  wire [1:0]        _GEN_443 = {{~_GEN_5}, {Register_inst2[89]}};
  wire [1:0]        _GEN_444 = {{~_GEN_5}, {Register_inst2[88]}};
  wire [1:0]        _GEN_445 = {{~_GEN_5}, {Register_inst2[87]}};
  wire [1:0]        _GEN_446 = {{~_GEN_5}, {Register_inst2[86]}};
  wire [1:0]        _GEN_447 = {{~_GEN_5}, {Register_inst2[85]}};
  wire [1:0]        _GEN_448 = {{~_GEN_5}, {Register_inst2[84]}};
  wire [1:0]        _GEN_449 = {{~_GEN_5}, {Register_inst2[83]}};
  wire [1:0]        _GEN_450 = {{~_GEN_5}, {Register_inst2[82]}};
  wire [1:0]        _GEN_451 = {{~_GEN_5}, {Register_inst2[81]}};
  wire [1:0]        _GEN_452 = {{~_GEN_5}, {Register_inst2[80]}};
  wire [1:0]        _GEN_453 = {{~_GEN_5}, {Register_inst2[79]}};
  wire [1:0]        _GEN_454 = {{~_GEN_5}, {Register_inst2[78]}};
  wire [1:0]        _GEN_455 = {{~_GEN_5}, {Register_inst2[77]}};
  wire [1:0]        _GEN_456 = {{~_GEN_5}, {Register_inst2[76]}};
  wire [1:0]        _GEN_457 = {{~_GEN_5}, {Register_inst2[75]}};
  wire [1:0]        _GEN_458 = {{~_GEN_5}, {Register_inst2[74]}};
  wire [1:0]        _GEN_459 = {{~_GEN_5}, {Register_inst2[73]}};
  wire [1:0]        _GEN_460 = {{~_GEN_5}, {Register_inst2[72]}};
  wire [1:0]        _GEN_461 = {{~_GEN_5}, {Register_inst2[71]}};
  wire [1:0]        _GEN_462 = {{~_GEN_5}, {Register_inst2[70]}};
  wire [1:0]        _GEN_463 = {{~_GEN_5}, {Register_inst2[69]}};
  wire [1:0]        _GEN_464 = {{~_GEN_5}, {Register_inst2[68]}};
  wire [1:0]        _GEN_465 = {{~_GEN_5}, {Register_inst2[67]}};
  wire [1:0]        _GEN_466 = {{~_GEN_5}, {Register_inst2[66]}};
  wire [1:0]        _GEN_467 = {{~_GEN_5}, {Register_inst2[65]}};
  wire [1:0]        _GEN_468 = {{~_GEN_5}, {Register_inst2[64]}};
  wire [1:0]        _GEN_469 = {{~_GEN_5}, {Register_inst2[63]}};
  wire [1:0]        _GEN_470 = {{~_GEN_5}, {Register_inst2[62]}};
  wire [1:0]        _GEN_471 = {{~_GEN_5}, {Register_inst2[61]}};
  wire [1:0]        _GEN_472 = {{~_GEN_5}, {Register_inst2[60]}};
  wire [1:0]        _GEN_473 = {{~_GEN_5}, {Register_inst2[59]}};
  wire [1:0]        _GEN_474 = {{~_GEN_5}, {Register_inst2[58]}};
  wire [1:0]        _GEN_475 = {{~_GEN_5}, {Register_inst2[57]}};
  wire [1:0]        _GEN_476 = {{~_GEN_5}, {Register_inst2[56]}};
  wire [1:0]        _GEN_477 = {{~_GEN_5}, {Register_inst2[55]}};
  wire [1:0]        _GEN_478 = {{~_GEN_5}, {Register_inst2[54]}};
  wire [1:0]        _GEN_479 = {{~_GEN_5}, {Register_inst2[53]}};
  wire [1:0]        _GEN_480 = {{~_GEN_5}, {Register_inst2[52]}};
  wire [1:0]        _GEN_481 = {{~_GEN_5}, {Register_inst2[51]}};
  wire [1:0]        _GEN_482 = {{~_GEN_5}, {Register_inst2[50]}};
  wire [1:0]        _GEN_483 = {{~_GEN_5}, {Register_inst2[49]}};
  wire [1:0]        _GEN_484 = {{~_GEN_5}, {Register_inst2[48]}};
  wire [1:0]        _GEN_485 = {{~_GEN_5}, {Register_inst2[47]}};
  wire [1:0]        _GEN_486 = {{~_GEN_5}, {Register_inst2[46]}};
  wire [1:0]        _GEN_487 = {{~_GEN_5}, {Register_inst2[45]}};
  wire [1:0]        _GEN_488 = {{~_GEN_5}, {Register_inst2[44]}};
  wire [1:0]        _GEN_489 = {{~_GEN_5}, {Register_inst2[43]}};
  wire [1:0]        _GEN_490 = {{~_GEN_5}, {Register_inst2[42]}};
  wire [1:0]        _GEN_491 = {{~_GEN_5}, {Register_inst2[41]}};
  wire [1:0]        _GEN_492 = {{~_GEN_5}, {Register_inst2[40]}};
  wire [1:0]        _GEN_493 = {{~_GEN_5}, {Register_inst2[39]}};
  wire [1:0]        _GEN_494 = {{~_GEN_5}, {Register_inst2[38]}};
  wire [1:0]        _GEN_495 = {{~_GEN_5}, {Register_inst2[37]}};
  wire [1:0]        _GEN_496 = {{~_GEN_5}, {Register_inst2[36]}};
  wire [1:0]        _GEN_497 = {{~_GEN_5}, {Register_inst2[35]}};
  wire [1:0]        _GEN_498 = {{~_GEN_5}, {Register_inst2[34]}};
  wire [1:0]        _GEN_499 = {{~_GEN_5}, {Register_inst2[33]}};
  wire [1:0]        _GEN_500 = {{~_GEN_5}, {Register_inst2[32]}};
  wire [1:0]        _GEN_501 = {{~_GEN_5}, {Register_inst2[31]}};
  wire [1:0]        _GEN_502 = {{~_GEN_5}, {Register_inst2[30]}};
  wire [1:0]        _GEN_503 = {{~_GEN_5}, {Register_inst2[29]}};
  wire [1:0]        _GEN_504 = {{~_GEN_5}, {Register_inst2[28]}};
  wire [1:0]        _GEN_505 = {{~_GEN_5}, {Register_inst2[27]}};
  wire [1:0]        _GEN_506 = {{~_GEN_5}, {Register_inst2[26]}};
  wire [1:0]        _GEN_507 = {{~_GEN_5}, {Register_inst2[25]}};
  wire [1:0]        _GEN_508 = {{~_GEN_5}, {Register_inst2[24]}};
  wire [1:0]        _GEN_509 = {{~_GEN_5}, {Register_inst2[23]}};
  wire [1:0]        _GEN_510 = {{~_GEN_5}, {Register_inst2[22]}};
  wire [1:0]        _GEN_511 = {{~_GEN_5}, {Register_inst2[21]}};
  wire [1:0]        _GEN_512 = {{~_GEN_5}, {Register_inst2[20]}};
  wire [1:0]        _GEN_513 = {{~_GEN_5}, {Register_inst2[19]}};
  wire [1:0]        _GEN_514 = {{~_GEN_5}, {Register_inst2[18]}};
  wire [1:0]        _GEN_515 = {{~_GEN_5}, {Register_inst2[17]}};
  wire [1:0]        _GEN_516 = {{~_GEN_5}, {Register_inst2[16]}};
  wire [1:0]        _GEN_517 = {{~_GEN_5}, {Register_inst2[15]}};
  wire [1:0]        _GEN_518 = {{~_GEN_5}, {Register_inst2[14]}};
  wire [1:0]        _GEN_519 = {{~_GEN_5}, {Register_inst2[13]}};
  wire [1:0]        _GEN_520 = {{~_GEN_5}, {Register_inst2[12]}};
  wire [1:0]        _GEN_521 = {{~_GEN_5}, {Register_inst2[11]}};
  wire [1:0]        _GEN_522 = {{~_GEN_5}, {Register_inst2[10]}};
  wire [1:0]        _GEN_523 = {{~_GEN_5}, {Register_inst2[9]}};
  wire [1:0]        _GEN_524 = {{~_GEN_5}, {Register_inst2[8]}};
  wire [1:0]        _GEN_525 = {{~_GEN_5}, {Register_inst2[7]}};
  wire [1:0]        _GEN_526 = {{~_GEN_5}, {Register_inst2[6]}};
  wire [1:0]        _GEN_527 = {{~_GEN_5}, {Register_inst2[5]}};
  wire [1:0]        _GEN_528 = {{~_GEN_5}, {Register_inst2[4]}};
  wire [1:0]        _GEN_529 = {{~_GEN_5}, {Register_inst2[3]}};
  wire [1:0]        _GEN_530 = {{~_GEN_5}, {Register_inst2[2]}};
  wire [1:0]        _GEN_531 = {{~_GEN_5}, {Register_inst2[1]}};
  wire [1:0]        _GEN_532 = {{~_GEN_5}, {Register_inst2[0]}};
  wire [255:0]      _GEN_533 =
    {_GEN_277[&(Register_inst3[11:4])],
     _GEN_278[Register_inst3[11:4] == 8'hFE],
     _GEN_279[Register_inst3[11:4] == 8'hFD],
     _GEN_280[Register_inst3[11:4] == 8'hFC],
     _GEN_281[Register_inst3[11:4] == 8'hFB],
     _GEN_282[Register_inst3[11:4] == 8'hFA],
     _GEN_283[Register_inst3[11:4] == 8'hF9],
     _GEN_284[Register_inst3[11:4] == 8'hF8],
     _GEN_285[Register_inst3[11:4] == 8'hF7],
     _GEN_286[Register_inst3[11:4] == 8'hF6],
     _GEN_287[Register_inst3[11:4] == 8'hF5],
     _GEN_288[Register_inst3[11:4] == 8'hF4],
     _GEN_289[Register_inst3[11:4] == 8'hF3],
     _GEN_290[Register_inst3[11:4] == 8'hF2],
     _GEN_291[Register_inst3[11:4] == 8'hF1],
     _GEN_292[Register_inst3[11:4] == 8'hF0],
     _GEN_293[Register_inst3[11:4] == 8'hEF],
     _GEN_294[Register_inst3[11:4] == 8'hEE],
     _GEN_295[Register_inst3[11:4] == 8'hED],
     _GEN_296[Register_inst3[11:4] == 8'hEC],
     _GEN_297[Register_inst3[11:4] == 8'hEB],
     _GEN_298[Register_inst3[11:4] == 8'hEA],
     _GEN_299[Register_inst3[11:4] == 8'hE9],
     _GEN_300[Register_inst3[11:4] == 8'hE8],
     _GEN_301[Register_inst3[11:4] == 8'hE7],
     _GEN_302[Register_inst3[11:4] == 8'hE6],
     _GEN_303[Register_inst3[11:4] == 8'hE5],
     _GEN_304[Register_inst3[11:4] == 8'hE4],
     _GEN_305[Register_inst3[11:4] == 8'hE3],
     _GEN_306[Register_inst3[11:4] == 8'hE2],
     _GEN_307[Register_inst3[11:4] == 8'hE1],
     _GEN_308[Register_inst3[11:4] == 8'hE0],
     _GEN_309[Register_inst3[11:4] == 8'hDF],
     _GEN_310[Register_inst3[11:4] == 8'hDE],
     _GEN_311[Register_inst3[11:4] == 8'hDD],
     _GEN_312[Register_inst3[11:4] == 8'hDC],
     _GEN_313[Register_inst3[11:4] == 8'hDB],
     _GEN_314[Register_inst3[11:4] == 8'hDA],
     _GEN_315[Register_inst3[11:4] == 8'hD9],
     _GEN_316[Register_inst3[11:4] == 8'hD8],
     _GEN_317[Register_inst3[11:4] == 8'hD7],
     _GEN_318[Register_inst3[11:4] == 8'hD6],
     _GEN_319[Register_inst3[11:4] == 8'hD5],
     _GEN_320[Register_inst3[11:4] == 8'hD4],
     _GEN_321[Register_inst3[11:4] == 8'hD3],
     _GEN_322[Register_inst3[11:4] == 8'hD2],
     _GEN_323[Register_inst3[11:4] == 8'hD1],
     _GEN_324[Register_inst3[11:4] == 8'hD0],
     _GEN_325[Register_inst3[11:4] == 8'hCF],
     _GEN_326[Register_inst3[11:4] == 8'hCE],
     _GEN_327[Register_inst3[11:4] == 8'hCD],
     _GEN_328[Register_inst3[11:4] == 8'hCC],
     _GEN_329[Register_inst3[11:4] == 8'hCB],
     _GEN_330[Register_inst3[11:4] == 8'hCA],
     _GEN_331[Register_inst3[11:4] == 8'hC9],
     _GEN_332[Register_inst3[11:4] == 8'hC8],
     _GEN_333[Register_inst3[11:4] == 8'hC7],
     _GEN_334[Register_inst3[11:4] == 8'hC6],
     _GEN_335[Register_inst3[11:4] == 8'hC5],
     _GEN_336[Register_inst3[11:4] == 8'hC4],
     _GEN_337[Register_inst3[11:4] == 8'hC3],
     _GEN_338[Register_inst3[11:4] == 8'hC2],
     _GEN_339[Register_inst3[11:4] == 8'hC1],
     _GEN_340[Register_inst3[11:4] == 8'hC0],
     _GEN_341[Register_inst3[11:4] == 8'hBF],
     _GEN_342[Register_inst3[11:4] == 8'hBE],
     _GEN_343[Register_inst3[11:4] == 8'hBD],
     _GEN_344[Register_inst3[11:4] == 8'hBC],
     _GEN_345[Register_inst3[11:4] == 8'hBB],
     _GEN_346[Register_inst3[11:4] == 8'hBA],
     _GEN_347[Register_inst3[11:4] == 8'hB9],
     _GEN_348[Register_inst3[11:4] == 8'hB8],
     _GEN_349[Register_inst3[11:4] == 8'hB7],
     _GEN_350[Register_inst3[11:4] == 8'hB6],
     _GEN_351[Register_inst3[11:4] == 8'hB5],
     _GEN_352[Register_inst3[11:4] == 8'hB4],
     _GEN_353[Register_inst3[11:4] == 8'hB3],
     _GEN_354[Register_inst3[11:4] == 8'hB2],
     _GEN_355[Register_inst3[11:4] == 8'hB1],
     _GEN_356[Register_inst3[11:4] == 8'hB0],
     _GEN_357[Register_inst3[11:4] == 8'hAF],
     _GEN_358[Register_inst3[11:4] == 8'hAE],
     _GEN_359[Register_inst3[11:4] == 8'hAD],
     _GEN_360[Register_inst3[11:4] == 8'hAC],
     _GEN_361[Register_inst3[11:4] == 8'hAB],
     _GEN_362[Register_inst3[11:4] == 8'hAA],
     _GEN_363[Register_inst3[11:4] == 8'hA9],
     _GEN_364[Register_inst3[11:4] == 8'hA8],
     _GEN_365[Register_inst3[11:4] == 8'hA7],
     _GEN_366[Register_inst3[11:4] == 8'hA6],
     _GEN_367[Register_inst3[11:4] == 8'hA5],
     _GEN_368[Register_inst3[11:4] == 8'hA4],
     _GEN_369[Register_inst3[11:4] == 8'hA3],
     _GEN_370[Register_inst3[11:4] == 8'hA2],
     _GEN_371[Register_inst3[11:4] == 8'hA1],
     _GEN_372[Register_inst3[11:4] == 8'hA0],
     _GEN_373[Register_inst3[11:4] == 8'h9F],
     _GEN_374[Register_inst3[11:4] == 8'h9E],
     _GEN_375[Register_inst3[11:4] == 8'h9D],
     _GEN_376[Register_inst3[11:4] == 8'h9C],
     _GEN_377[Register_inst3[11:4] == 8'h9B],
     _GEN_378[Register_inst3[11:4] == 8'h9A],
     _GEN_379[Register_inst3[11:4] == 8'h99],
     _GEN_380[Register_inst3[11:4] == 8'h98],
     _GEN_381[Register_inst3[11:4] == 8'h97],
     _GEN_382[Register_inst3[11:4] == 8'h96],
     _GEN_383[Register_inst3[11:4] == 8'h95],
     _GEN_384[Register_inst3[11:4] == 8'h94],
     _GEN_385[Register_inst3[11:4] == 8'h93],
     _GEN_386[Register_inst3[11:4] == 8'h92],
     _GEN_387[Register_inst3[11:4] == 8'h91],
     _GEN_388[Register_inst3[11:4] == 8'h90],
     _GEN_389[Register_inst3[11:4] == 8'h8F],
     _GEN_390[Register_inst3[11:4] == 8'h8E],
     _GEN_391[Register_inst3[11:4] == 8'h8D],
     _GEN_392[Register_inst3[11:4] == 8'h8C],
     _GEN_393[Register_inst3[11:4] == 8'h8B],
     _GEN_394[Register_inst3[11:4] == 8'h8A],
     _GEN_395[Register_inst3[11:4] == 8'h89],
     _GEN_396[Register_inst3[11:4] == 8'h88],
     _GEN_397[Register_inst3[11:4] == 8'h87],
     _GEN_398[Register_inst3[11:4] == 8'h86],
     _GEN_399[Register_inst3[11:4] == 8'h85],
     _GEN_400[Register_inst3[11:4] == 8'h84],
     _GEN_401[Register_inst3[11:4] == 8'h83],
     _GEN_402[Register_inst3[11:4] == 8'h82],
     _GEN_403[Register_inst3[11:4] == 8'h81],
     _GEN_404[Register_inst3[11:4] == 8'h80],
     _GEN_405[Register_inst3[11:4] == 8'h7F],
     _GEN_406[Register_inst3[11:4] == 8'h7E],
     _GEN_407[Register_inst3[11:4] == 8'h7D],
     _GEN_408[Register_inst3[11:4] == 8'h7C],
     _GEN_409[Register_inst3[11:4] == 8'h7B],
     _GEN_410[Register_inst3[11:4] == 8'h7A],
     _GEN_411[Register_inst3[11:4] == 8'h79],
     _GEN_412[Register_inst3[11:4] == 8'h78],
     _GEN_413[Register_inst3[11:4] == 8'h77],
     _GEN_414[Register_inst3[11:4] == 8'h76],
     _GEN_415[Register_inst3[11:4] == 8'h75],
     _GEN_416[Register_inst3[11:4] == 8'h74],
     _GEN_417[Register_inst3[11:4] == 8'h73],
     _GEN_418[Register_inst3[11:4] == 8'h72],
     _GEN_419[Register_inst3[11:4] == 8'h71],
     _GEN_420[Register_inst3[11:4] == 8'h70],
     _GEN_421[Register_inst3[11:4] == 8'h6F],
     _GEN_422[Register_inst3[11:4] == 8'h6E],
     _GEN_423[Register_inst3[11:4] == 8'h6D],
     _GEN_424[Register_inst3[11:4] == 8'h6C],
     _GEN_425[Register_inst3[11:4] == 8'h6B],
     _GEN_426[Register_inst3[11:4] == 8'h6A],
     _GEN_427[Register_inst3[11:4] == 8'h69],
     _GEN_428[Register_inst3[11:4] == 8'h68],
     _GEN_429[Register_inst3[11:4] == 8'h67],
     _GEN_430[Register_inst3[11:4] == 8'h66],
     _GEN_431[Register_inst3[11:4] == 8'h65],
     _GEN_432[Register_inst3[11:4] == 8'h64],
     _GEN_433[Register_inst3[11:4] == 8'h63],
     _GEN_434[Register_inst3[11:4] == 8'h62],
     _GEN_435[Register_inst3[11:4] == 8'h61],
     _GEN_436[Register_inst3[11:4] == 8'h60],
     _GEN_437[Register_inst3[11:4] == 8'h5F],
     _GEN_438[Register_inst3[11:4] == 8'h5E],
     _GEN_439[Register_inst3[11:4] == 8'h5D],
     _GEN_440[Register_inst3[11:4] == 8'h5C],
     _GEN_441[Register_inst3[11:4] == 8'h5B],
     _GEN_442[Register_inst3[11:4] == 8'h5A],
     _GEN_443[Register_inst3[11:4] == 8'h59],
     _GEN_444[Register_inst3[11:4] == 8'h58],
     _GEN_445[Register_inst3[11:4] == 8'h57],
     _GEN_446[Register_inst3[11:4] == 8'h56],
     _GEN_447[Register_inst3[11:4] == 8'h55],
     _GEN_448[Register_inst3[11:4] == 8'h54],
     _GEN_449[Register_inst3[11:4] == 8'h53],
     _GEN_450[Register_inst3[11:4] == 8'h52],
     _GEN_451[Register_inst3[11:4] == 8'h51],
     _GEN_452[Register_inst3[11:4] == 8'h50],
     _GEN_453[Register_inst3[11:4] == 8'h4F],
     _GEN_454[Register_inst3[11:4] == 8'h4E],
     _GEN_455[Register_inst3[11:4] == 8'h4D],
     _GEN_456[Register_inst3[11:4] == 8'h4C],
     _GEN_457[Register_inst3[11:4] == 8'h4B],
     _GEN_458[Register_inst3[11:4] == 8'h4A],
     _GEN_459[Register_inst3[11:4] == 8'h49],
     _GEN_460[Register_inst3[11:4] == 8'h48],
     _GEN_461[Register_inst3[11:4] == 8'h47],
     _GEN_462[Register_inst3[11:4] == 8'h46],
     _GEN_463[Register_inst3[11:4] == 8'h45],
     _GEN_464[Register_inst3[11:4] == 8'h44],
     _GEN_465[Register_inst3[11:4] == 8'h43],
     _GEN_466[Register_inst3[11:4] == 8'h42],
     _GEN_467[Register_inst3[11:4] == 8'h41],
     _GEN_468[Register_inst3[11:4] == 8'h40],
     _GEN_469[Register_inst3[11:4] == 8'h3F],
     _GEN_470[Register_inst3[11:4] == 8'h3E],
     _GEN_471[Register_inst3[11:4] == 8'h3D],
     _GEN_472[Register_inst3[11:4] == 8'h3C],
     _GEN_473[Register_inst3[11:4] == 8'h3B],
     _GEN_474[Register_inst3[11:4] == 8'h3A],
     _GEN_475[Register_inst3[11:4] == 8'h39],
     _GEN_476[Register_inst3[11:4] == 8'h38],
     _GEN_477[Register_inst3[11:4] == 8'h37],
     _GEN_478[Register_inst3[11:4] == 8'h36],
     _GEN_479[Register_inst3[11:4] == 8'h35],
     _GEN_480[Register_inst3[11:4] == 8'h34],
     _GEN_481[Register_inst3[11:4] == 8'h33],
     _GEN_482[Register_inst3[11:4] == 8'h32],
     _GEN_483[Register_inst3[11:4] == 8'h31],
     _GEN_484[Register_inst3[11:4] == 8'h30],
     _GEN_485[Register_inst3[11:4] == 8'h2F],
     _GEN_486[Register_inst3[11:4] == 8'h2E],
     _GEN_487[Register_inst3[11:4] == 8'h2D],
     _GEN_488[Register_inst3[11:4] == 8'h2C],
     _GEN_489[Register_inst3[11:4] == 8'h2B],
     _GEN_490[Register_inst3[11:4] == 8'h2A],
     _GEN_491[Register_inst3[11:4] == 8'h29],
     _GEN_492[Register_inst3[11:4] == 8'h28],
     _GEN_493[Register_inst3[11:4] == 8'h27],
     _GEN_494[Register_inst3[11:4] == 8'h26],
     _GEN_495[Register_inst3[11:4] == 8'h25],
     _GEN_496[Register_inst3[11:4] == 8'h24],
     _GEN_497[Register_inst3[11:4] == 8'h23],
     _GEN_498[Register_inst3[11:4] == 8'h22],
     _GEN_499[Register_inst3[11:4] == 8'h21],
     _GEN_500[Register_inst3[11:4] == 8'h20],
     _GEN_501[Register_inst3[11:4] == 8'h1F],
     _GEN_502[Register_inst3[11:4] == 8'h1E],
     _GEN_503[Register_inst3[11:4] == 8'h1D],
     _GEN_504[Register_inst3[11:4] == 8'h1C],
     _GEN_505[Register_inst3[11:4] == 8'h1B],
     _GEN_506[Register_inst3[11:4] == 8'h1A],
     _GEN_507[Register_inst3[11:4] == 8'h19],
     _GEN_508[Register_inst3[11:4] == 8'h18],
     _GEN_509[Register_inst3[11:4] == 8'h17],
     _GEN_510[Register_inst3[11:4] == 8'h16],
     _GEN_511[Register_inst3[11:4] == 8'h15],
     _GEN_512[Register_inst3[11:4] == 8'h14],
     _GEN_513[Register_inst3[11:4] == 8'h13],
     _GEN_514[Register_inst3[11:4] == 8'h12],
     _GEN_515[Register_inst3[11:4] == 8'h11],
     _GEN_516[Register_inst3[11:4] == 8'h10],
     _GEN_517[Register_inst3[11:4] == 8'hF],
     _GEN_518[Register_inst3[11:4] == 8'hE],
     _GEN_519[Register_inst3[11:4] == 8'hD],
     _GEN_520[Register_inst3[11:4] == 8'hC],
     _GEN_521[Register_inst3[11:4] == 8'hB],
     _GEN_522[Register_inst3[11:4] == 8'hA],
     _GEN_523[Register_inst3[11:4] == 8'h9],
     _GEN_524[Register_inst3[11:4] == 8'h8],
     _GEN_525[Register_inst3[11:4] == 8'h7],
     _GEN_526[Register_inst3[11:4] == 8'h6],
     _GEN_527[Register_inst3[11:4] == 8'h5],
     _GEN_528[Register_inst3[11:4] == 8'h4],
     _GEN_529[Register_inst3[11:4] == 8'h3],
     _GEN_530[Register_inst3[11:4] == 8'h2],
     _GEN_531[Register_inst3[11:4] == 8'h1],
     _GEN_532[Register_inst3[11:4] == 8'h0]};
  wire [1:0][63:0]  _GEN_534 = {{nasti_r_data.data}, {Register_inst6[1'h1]}};
  wire [1:0][63:0]  _GEN_535 = {{nasti_r_data.data}, {Register_inst6[1'h0]}};
  always_ff @(posedge CLK) begin
    if (_GEN_15)
      Register_inst3 <= cpu_req.data.addr;
    Register_inst7 <= _GEN_5;
    if (_GEN_6) begin
      Register_inst1 <= _GEN_276;
      Register_inst2 <= _GEN_533;
    end
    if (_GEN_15)
      Register_inst5 <= cpu_req.data.mask;
    if (_GEN_4 & nasti_r_valid)
      Register_inst6 <= {{_GEN_534[_Counter_inst0_O]}, {_GEN_535[~_Counter_inst0_O]}};
    if (_GEN_15)
      Register_inst4 <= cpu_req.data.data;
    Register_inst8 <= _GEN_9;
    if (Register_inst8)
      Register_inst9 <=
        {_ArrayMaskMem_inst3_RDATA,
         _ArrayMaskMem_inst2_RDATA,
         _ArrayMaskMem_inst1_RDATA,
         _ArrayMaskMem_inst0_RDATA};
  end // always_ff @(posedge)
  initial begin
    Register_inst3 = 32'h0;
    Register_inst7 = 1'h0;
    Register_inst1 = 256'h0;
    Register_inst2 = 256'h0;
    Register_inst5 = 4'h0;
    Register_inst0 = 3'h0;
    Register_inst6 = {64'h0, 64'h0};
    Register_inst4 = 32'h0;
    Register_inst8 = 1'h0;
    Register_inst9 =
      {8'h0,
       8'h0,
       8'h0,
       8'h0,
       8'h0,
       8'h0,
       8'h0,
       8'h0,
       8'h0,
       8'h0,
       8'h0,
       8'h0,
       8'h0,
       8'h0,
       8'h0,
       8'h0};
  end // initial
  wire [1:0][7:0]   _GEN_536 =
    {{_ArrayMaskMem_inst0_RDATA[2'h0]}, {Register_inst9[4'h0]}};
  wire [1:0][7:0]   _GEN_537 =
    {{_ArrayMaskMem_inst0_RDATA[2'h1]}, {Register_inst9[4'h1]}};
  wire [1:0][7:0]   _GEN_538 =
    {{_ArrayMaskMem_inst0_RDATA[2'h2]}, {Register_inst9[4'h2]}};
  wire [1:0][7:0]   _GEN_539 =
    {{_ArrayMaskMem_inst0_RDATA[2'h3]}, {Register_inst9[4'h3]}};
  wire [1:0][7:0]   _GEN_540 =
    {{_ArrayMaskMem_inst1_RDATA[2'h0]}, {Register_inst9[4'h4]}};
  wire [1:0][7:0]   _GEN_541 =
    {{_ArrayMaskMem_inst1_RDATA[2'h1]}, {Register_inst9[4'h5]}};
  wire [1:0][7:0]   _GEN_542 =
    {{_ArrayMaskMem_inst1_RDATA[2'h2]}, {Register_inst9[4'h6]}};
  wire [1:0][7:0]   _GEN_543 =
    {{_ArrayMaskMem_inst1_RDATA[2'h3]}, {Register_inst9[4'h7]}};
  wire [1:0][7:0]   _GEN_544 =
    {{_ArrayMaskMem_inst2_RDATA[2'h0]}, {Register_inst9[4'h8]}};
  wire [1:0][7:0]   _GEN_545 =
    {{_ArrayMaskMem_inst2_RDATA[2'h1]}, {Register_inst9[4'h9]}};
  wire [1:0][7:0]   _GEN_546 =
    {{_ArrayMaskMem_inst2_RDATA[2'h2]}, {Register_inst9[4'hA]}};
  wire [1:0][7:0]   _GEN_547 =
    {{_ArrayMaskMem_inst2_RDATA[2'h3]}, {Register_inst9[4'hB]}};
  wire [1:0][7:0]   _GEN_548 =
    {{_ArrayMaskMem_inst3_RDATA[2'h0]}, {Register_inst9[4'hC]}};
  wire [1:0][7:0]   _GEN_549 =
    {{_ArrayMaskMem_inst3_RDATA[2'h1]}, {Register_inst9[4'hD]}};
  wire [1:0][7:0]   _GEN_550 =
    {{_ArrayMaskMem_inst3_RDATA[2'h2]}, {Register_inst9[4'hE]}};
  wire [1:0][7:0]   _GEN_551 =
    {{_ArrayMaskMem_inst3_RDATA[2'h3]}, {Register_inst9[4'hF]}};
  wire [127:0]      _GEN_552 = /*cast(bit[127:0])*/Register_inst6;
  wire [1:0][127:0] _GEN_553 =
    {{_GEN_552},
     {{_GEN_551[Register_inst8],
       _GEN_550[Register_inst8],
       _GEN_549[Register_inst8],
       _GEN_548[Register_inst8],
       _GEN_547[Register_inst8],
       _GEN_546[Register_inst8],
       _GEN_545[Register_inst8],
       _GEN_544[Register_inst8],
       _GEN_543[Register_inst8],
       _GEN_542[Register_inst8],
       _GEN_541[Register_inst8],
       _GEN_540[Register_inst8],
       _GEN_539[Register_inst8],
       _GEN_538[Register_inst8],
       _GEN_537[Register_inst8],
       _GEN_536[Register_inst8]}}};
  wire [127:0]      _GEN_554 = _GEN_553[Register_inst7];
  wire [3:0][31:0]  _GEN_555 =
    {{_GEN_554[127:96]}, {_GEN_554[95:64]}, {_GEN_554[63:32]}, {_GEN_554[31:0]}};
  wire struct packed {logic [31:0] data; } _GEN_556;
  assign _GEN_556.data = _GEN_555[Register_inst3[3:2]];
  wire struct packed {logic valid; struct packed {logic [31:0] data; } data; } _GEN_557;
  assign _GEN_557.valid = _GEN_15;
  assign _GEN_557.data = _GEN_556;
  wire
    struct packed {logic [4:0] id; logic user; logic [31:0] addr; logic [7:0] length; logic [2:0] size; logic [1:0] burst; logic lock; logic [3:0] cache; logic [2:0] prot; logic [3:0] qos; logic [3:0] region; }
    _GEN_558;
  assign _GEN_558.id = 5'h0;
  assign _GEN_558.user = 1'h0;
  assign _GEN_558.addr = {_Memory_inst0_RDATA.tag, Register_inst3[11:4], 4'h0};
  assign _GEN_558.length = 8'h1;
  assign _GEN_558.size = 3'h3;
  assign _GEN_558.burst = 2'h1;
  assign _GEN_558.lock = 1'h0;
  assign _GEN_558.cache = 4'h0;
  assign _GEN_558.prot = 3'h0;
  assign _GEN_558.qos = 4'h0;
  assign _GEN_558.region = 4'h0;
  wire [1:0][63:0]  _GEN_559 = {{_GEN_554[127:64]}, {_GEN_554[63:0]}};
  wire
    struct packed {logic [4:0] id; logic [7:0] strb; logic user; logic [63:0] data; logic last; }
    _GEN_560;
  assign _GEN_560.id = 5'h0;
  assign _GEN_560.strb = 8'hFF;
  assign _GEN_560.user = 1'h0;
  assign _GEN_560.data = _GEN_559[_Counter_inst1_O];
  assign _GEN_560.last = _Counter_inst1_COUT;
  wire
    struct packed {logic [4:0] id; logic user; logic [31:0] addr; logic [7:0] length; logic [2:0] size; logic [1:0] burst; logic lock; logic [3:0] cache; logic [2:0] prot; logic [3:0] qos; logic [3:0] region; }
    _GEN_561;
  assign _GEN_561.id = 5'h0;
  assign _GEN_561.user = 1'h0;
  assign _GEN_561.addr = {Register_inst3[31:4], 4'h0};
  assign _GEN_561.length = 8'h1;
  assign _GEN_561.size = 3'h3;
  assign _GEN_561.burst = 2'h1;
  assign _GEN_561.lock = 1'h0;
  assign _GEN_561.cache = 4'h0;
  assign _GEN_561.prot = 3'h0;
  assign _GEN_561.qos = 4'h0;
  assign _GEN_561.region = 4'h0;
  always @(posedge CLK) begin
      $display("resp.valid=%x", _GEN_15);
  end
  always @(posedge CLK) begin
      $display("[%0t]: valid = %x", $time, _GEN_15);
  end
  always @(posedge CLK) begin
      $display("[%0t]: is_idle = %x, is_read = %x, hit = %x, is_alloc_reg = %x, ~cpu_mask.O.reduce_or() = %x", $time, _GEN, _GEN_8, hit, Register_inst7, Register_inst5 == 4'h0);
  end
  always @(posedge CLK) begin
      if (_GEN_15 & Register_inst7) $display("[%0t]: refill_buf.O=%x, %x", $time, Register_inst6[1'h0], Register_inst6[1'h1]);
  end
  always @(posedge CLK) begin
      if (_GEN_15 & Register_inst7) $display("[%0t]: read=%x", $time, _GEN_554);
  end
  Counter Counter_inst0 (
    .CLK   (CLK),
    .CE    (_GEN_4 & nasti_r_valid),
    .RESET (RESET),
    .O     (_Counter_inst0_O),
    .COUT  (_Counter_inst0_COUT)
  );
  Memory Memory_inst0 (
    .RADDR (cpu_req.data.addr[11:4]),
    .CLK   (CLK),
    .RE    (_GEN_9),
    .WADDR (Register_inst3[11:4]),
    .WDATA (wmeta),
    .WE    (_GEN_6 & _GEN_5),
    .RDATA (_Memory_inst0_RDATA)
  );
  Counter Counter_inst1 (
    .CLK   (CLK),
    .CE    (nasti_w_ready & _GEN_1),
    .RESET (RESET),
    .O     (_Counter_inst1_O),
    .COUT  (_Counter_inst1_COUT)
  );
  ArrayMaskMem ArrayMaskMem_inst0 (
    .RADDR (cpu_req.data.addr[11:4]),
    .CLK   (CLK),
    .RE    (_GEN_9),
    .WADDR (Register_inst3[11:4]),
    .WDATA ({{_GEN_17[31:24]}, {_GEN_17[23:16]}, {_GEN_17[15:8]}, {_GEN_17[7:0]}}),
    .WMASK (_GEN_19[3:0]),
    .WE    (_GEN_6),
    .RDATA (_ArrayMaskMem_inst0_RDATA)
  );
  ArrayMaskMem ArrayMaskMem_inst1 (
    .RADDR (cpu_req.data.addr[11:4]),
    .CLK   (CLK),
    .RE    (_GEN_9),
    .WADDR (Register_inst3[11:4]),
    .WDATA ({{_GEN_17[63:56]}, {_GEN_17[55:48]}, {_GEN_17[47:40]}, {_GEN_17[39:32]}}),
    .WMASK (_GEN_19[7:4]),
    .WE    (_GEN_6),
    .RDATA (_ArrayMaskMem_inst1_RDATA)
  );
  ArrayMaskMem ArrayMaskMem_inst2 (
    .RADDR (cpu_req.data.addr[11:4]),
    .CLK   (CLK),
    .RE    (_GEN_9),
    .WADDR (Register_inst3[11:4]),
    .WDATA ({{_GEN_17[95:88]}, {_GEN_17[87:80]}, {_GEN_17[79:72]}, {_GEN_17[71:64]}}),
    .WMASK (_GEN_19[11:8]),
    .WE    (_GEN_6),
    .RDATA (_ArrayMaskMem_inst2_RDATA)
  );
  ArrayMaskMem ArrayMaskMem_inst3 (
    .RADDR (cpu_req.data.addr[11:4]),
    .CLK   (CLK),
    .RE    (_GEN_9),
    .WADDR (Register_inst3[11:4]),
    .WDATA
      ({{_GEN_17[127:120]}, {_GEN_17[119:112]}, {_GEN_17[111:104]}, {_GEN_17[103:96]}}),
    .WMASK (_GEN_19[15:12]),
    .WE    (_GEN_6),
    .RDATA (_ArrayMaskMem_inst3_RDATA)
  );
  assign cpu_resp = _GEN_557;
  assign nasti_aw_valid = aw_valid;
  assign nasti_aw_data = _GEN_558;
  assign nasti_w_valid = _GEN_1;
  assign nasti_w_data = _GEN_560;
  assign nasti_b_ready = b_ready;
  assign nasti_ar_valid = ar_valid;
  assign nasti_ar_data = _GEN_561;
  assign nasti_r_ready = _GEN_4;
endmodule

module MemArbiter(
  input                                                                                                                                                                                                                 icache_aw_valid,
  input  struct packed {logic [4:0] id; logic user; logic [31:0] addr; logic [7:0] length; logic [2:0] size; logic [1:0] burst; logic lock; logic [3:0] cache; logic [2:0] prot; logic [3:0] qos; logic [3:0] region; } icache_aw_data,
  input                                                                                                                                                                                                                 icache_w_valid,
  input  struct packed {logic [4:0] id; logic [7:0] strb; logic user; logic [63:0] data; logic last; }                                                                                                                  icache_w_data,
  input                                                                                                                                                                                                                 icache_b_ready,
                                                                                                                                                                                                                        icache_ar_valid,
  input  struct packed {logic [4:0] id; logic user; logic [31:0] addr; logic [7:0] length; logic [2:0] size; logic [1:0] burst; logic lock; logic [3:0] cache; logic [2:0] prot; logic [3:0] qos; logic [3:0] region; } icache_ar_data,
  input                                                                                                                                                                                                                 icache_r_ready,
                                                                                                                                                                                                                        dcache_aw_valid,
  input  struct packed {logic [4:0] id; logic user; logic [31:0] addr; logic [7:0] length; logic [2:0] size; logic [1:0] burst; logic lock; logic [3:0] cache; logic [2:0] prot; logic [3:0] qos; logic [3:0] region; } dcache_aw_data,
  input                                                                                                                                                                                                                 dcache_w_valid,
  input  struct packed {logic [4:0] id; logic [7:0] strb; logic user; logic [63:0] data; logic last; }                                                                                                                  dcache_w_data,
  input                                                                                                                                                                                                                 dcache_b_ready,
                                                                                                                                                                                                                        dcache_ar_valid,
  input  struct packed {logic [4:0] id; logic user; logic [31:0] addr; logic [7:0] length; logic [2:0] size; logic [1:0] burst; logic lock; logic [3:0] cache; logic [2:0] prot; logic [3:0] qos; logic [3:0] region; } dcache_ar_data,
  input                                                                                                                                                                                                                 dcache_r_ready,
                                                                                                                                                                                                                        nasti_aw_ready,
                                                                                                                                                                                                                        nasti_w_ready,
                                                                                                                                                                                                                        nasti_b_valid,
  input  struct packed {logic [1:0] resp; logic [4:0] id; logic user; }                                                                                                                                                 nasti_b_data,
  input                                                                                                                                                                                                                 nasti_ar_ready,
                                                                                                                                                                                                                        nasti_r_valid,
  input  struct packed {logic [1:0] resp; logic [4:0] id; logic user; logic [63:0] data; logic last; }                                                                                                                  nasti_r_data,
  input                                                                                                                                                                                                                 CLK,
                                                                                                                                                                                                                        RESET,
  output                                                                                                                                                                                                                icache_aw_ready,
                                                                                                                                                                                                                        icache_w_ready,
                                                                                                                                                                                                                        icache_b_valid,
  output struct packed {logic [1:0] resp; logic [4:0] id; logic user; }                                                                                                                                                 icache_b_data,
  output                                                                                                                                                                                                                icache_ar_ready,
                                                                                                                                                                                                                        icache_r_valid,
  output struct packed {logic [1:0] resp; logic [4:0] id; logic user; logic [63:0] data; logic last; }                                                                                                                  icache_r_data,
  output                                                                                                                                                                                                                dcache_aw_ready,
                                                                                                                                                                                                                        dcache_w_ready,
                                                                                                                                                                                                                        dcache_b_valid,
  output struct packed {logic [1:0] resp; logic [4:0] id; logic user; }                                                                                                                                                 dcache_b_data,
  output                                                                                                                                                                                                                dcache_ar_ready,
                                                                                                                                                                                                                        dcache_r_valid,
  output struct packed {logic [1:0] resp; logic [4:0] id; logic user; logic [63:0] data; logic last; }                                                                                                                  dcache_r_data,
  output                                                                                                                                                                                                                nasti_aw_valid,
  output struct packed {logic [4:0] id; logic user; logic [31:0] addr; logic [7:0] length; logic [2:0] size; logic [1:0] burst; logic lock; logic [3:0] cache; logic [2:0] prot; logic [3:0] qos; logic [3:0] region; } nasti_aw_data,
  output                                                                                                                                                                                                                nasti_w_valid,
  output struct packed {logic [4:0] id; logic [7:0] strb; logic user; logic [63:0] data; logic last; }                                                                                                                  nasti_w_data,
  output                                                                                                                                                                                                                nasti_b_ready,
                                                                                                                                                                                                                        nasti_ar_valid,
  output struct packed {logic [4:0] id; logic user; logic [31:0] addr; logic [7:0] length; logic [2:0] size; logic [1:0] burst; logic lock; logic [3:0] cache; logic [2:0] prot; logic [3:0] qos; logic [3:0] region; } nasti_ar_data,
  output                                                                                                                                                                                                                nasti_r_ready
);

  wire             _GEN;
  wire             _GEN_0;
  reg  [2:0]       Register_inst0;
  wire struct packed {logic [1:0] resp; logic [4:0] id; logic user; } _GEN_1;
  assign _GEN_1.resp = 2'h0;
  assign _GEN_1.id = 5'h0;
  assign _GEN_1.user = 1'h0;
  wire             _GEN_2 = nasti_aw_ready & Register_inst0 == 3'h0;
  wire             _GEN_3 =
    icache_r_ready & Register_inst0 == 3'h1 | dcache_r_ready & Register_inst0 == 3'h2;
  wire             _GEN_4 = nasti_w_ready & Register_inst0 == 3'h3;
  wire             _GEN_5 = dcache_b_ready & Register_inst0 == 3'h4;
  reg  [2:0]       _GEN_6;
  always_comb begin
    _GEN_6 = Register_inst0;
    if (Register_inst0 == 3'h0) begin
      if (dcache_aw_valid & _GEN_2)
        _GEN_6 = 3'h3;
      else if (dcache_ar_valid & _GEN_0)
        _GEN_6 = 3'h2;
      else if (icache_ar_valid & _GEN)
        _GEN_6 = 3'h1;
    end
    else if (Register_inst0 == 3'h1) begin
      if (_GEN_3 & nasti_r_valid & nasti_r_data.last)
        _GEN_6 = 3'h0;
    end
    else if (Register_inst0 == 3'h2) begin
      if (_GEN_3 & nasti_r_valid & nasti_r_data.last)
        _GEN_6 = 3'h0;
    end
    else if (Register_inst0 == 3'h3) begin
      if (dcache_w_valid & _GEN_4 & dcache_w_data.last)
        _GEN_6 = 3'h4;
    end
    else if (Register_inst0 == 3'h4) begin
      if (_GEN_5 & nasti_b_valid)
        _GEN_6 = 3'h0;
    end
  end // always_comb
  always_ff @(posedge CLK)
    Register_inst0 <= _GEN_6;
  initial
    Register_inst0 = 3'h0;
  wire             _GEN_7 = dcache_aw_valid & Register_inst0 == 3'h0;
  assign _GEN_0 = nasti_ar_ready & ~_GEN_7 & Register_inst0 == 3'h0;
  assign _GEN = _GEN_0 & ~dcache_ar_valid;
  wire [1:0][4:0]  _GEN_8 = {{dcache_ar_data.id}, {icache_ar_data.id}};
  wire [1:0][31:0] _GEN_9 = {{dcache_ar_data.addr}, {icache_ar_data.addr}};
  wire [1:0][7:0]  _GEN_10 = {{dcache_ar_data.length}, {icache_ar_data.length}};
  wire [1:0][2:0]  _GEN_11 = {{dcache_ar_data.size}, {icache_ar_data.size}};
  wire
    struct packed {logic [4:0] id; logic user; logic [31:0] addr; logic [7:0] length; logic [2:0] size; logic [1:0] burst; logic lock; logic [3:0] cache; logic [2:0] prot; logic [3:0] qos; logic [3:0] region; }
    _GEN_12;
  assign _GEN_12.id = _GEN_8[dcache_ar_valid];
  assign _GEN_12.user = 1'h0;
  assign _GEN_12.addr = _GEN_9[dcache_ar_valid];
  assign _GEN_12.length = _GEN_10[dcache_ar_valid];
  assign _GEN_12.size = _GEN_11[dcache_ar_valid];
  assign _GEN_12.burst = 2'h1;
  assign _GEN_12.lock = 1'h0;
  assign _GEN_12.cache = 4'h0;
  assign _GEN_12.prot = 3'h0;
  assign _GEN_12.qos = 4'h0;
  assign _GEN_12.region = 4'h0;
  assign icache_aw_ready = 1'h0;
  assign icache_w_ready = 1'h0;
  assign icache_b_valid = 1'h0;
  assign icache_b_data = _GEN_1;
  assign icache_ar_ready = _GEN;
  assign icache_r_valid = nasti_r_valid & Register_inst0 == 3'h1;
  assign icache_r_data = nasti_r_data;
  assign dcache_aw_ready = _GEN_2;
  assign dcache_w_ready = _GEN_4;
  assign dcache_b_valid = nasti_b_valid & Register_inst0 == 3'h4;
  assign dcache_b_data = nasti_b_data;
  assign dcache_ar_ready = _GEN_0;
  assign dcache_r_valid = nasti_r_valid & Register_inst0 == 3'h2;
  assign dcache_r_data = nasti_r_data;
  assign nasti_aw_valid = _GEN_7;
  assign nasti_aw_data = dcache_aw_data;
  assign nasti_w_valid = dcache_w_valid & Register_inst0 == 3'h3;
  assign nasti_w_data = dcache_w_data;
  assign nasti_b_ready = _GEN_5;
  assign nasti_ar_valid =
    (icache_ar_valid | dcache_ar_valid) & ~_GEN_7 & Register_inst0 == 3'h0;
  assign nasti_ar_data = _GEN_12;
  assign nasti_r_ready = _GEN_3;
endmodule

module Tile(
  input  struct packed {logic valid; logic [31:0] data; }                                                                                                                                                               host_fromhost,
  input                                                                                                                                                                                                                 nasti_aw_ready,
                                                                                                                                                                                                                        nasti_w_ready,
                                                                                                                                                                                                                        nasti_b_valid,
  input  struct packed {logic [1:0] resp; logic [4:0] id; logic user; }                                                                                                                                                 nasti_b_data,
  input                                                                                                                                                                                                                 nasti_ar_ready,
                                                                                                                                                                                                                        nasti_r_valid,
  input  struct packed {logic [1:0] resp; logic [4:0] id; logic user; logic [63:0] data; logic last; }                                                                                                                  nasti_r_data,
  input                                                                                                                                                                                                                 CLK,
                                                                                                                                                                                                                        RESET,
  output [31:0]                                                                                                                                                                                                         host_tohost,
  output                                                                                                                                                                                                                nasti_aw_valid,
  output struct packed {logic [4:0] id; logic user; logic [31:0] addr; logic [7:0] length; logic [2:0] size; logic [1:0] burst; logic lock; logic [3:0] cache; logic [2:0] prot; logic [3:0] qos; logic [3:0] region; } nasti_aw_data,
  output                                                                                                                                                                                                                nasti_w_valid,
  output struct packed {logic [4:0] id; logic [7:0] strb; logic user; logic [63:0] data; logic last; }                                                                                                                  nasti_w_data,
  output                                                                                                                                                                                                                nasti_b_ready,
                                                                                                                                                                                                                        nasti_ar_valid,
  output struct packed {logic [4:0] id; logic user; logic [31:0] addr; logic [7:0] length; logic [2:0] size; logic [1:0] burst; logic lock; logic [3:0] cache; logic [2:0] prot; logic [3:0] qos; logic [3:0] region; } nasti_ar_data,
  output                                                                                                                                                                                                                nasti_r_ready
);

  wire _Core_inst0_icache_abort;
  wire
    struct packed {logic valid; struct packed {logic [31:0] addr; logic [31:0] data; logic [3:0] mask; } data; }
    _Core_inst0_icache_req;
  wire _Core_inst0_dcache_abort;
  wire
    struct packed {logic valid; struct packed {logic [31:0] addr; logic [31:0] data; logic [3:0] mask; } data; }
    _Core_inst0_dcache_req;
  wire struct packed {logic valid; struct packed {logic [31:0] data; } data; }
    _Cache_inst0_cpu_resp;
  wire _Cache_inst0_nasti_aw_valid;
  wire
    struct packed {logic [4:0] id; logic user; logic [31:0] addr; logic [7:0] length; logic [2:0] size; logic [1:0] burst; logic lock; logic [3:0] cache; logic [2:0] prot; logic [3:0] qos; logic [3:0] region; }
    _Cache_inst0_nasti_aw_data;
  wire _Cache_inst0_nasti_w_valid;
  wire
    struct packed {logic [4:0] id; logic [7:0] strb; logic user; logic [63:0] data; logic last; }
    _Cache_inst0_nasti_w_data;
  wire _Cache_inst0_nasti_b_ready;
  wire _Cache_inst0_nasti_ar_valid;
  wire
    struct packed {logic [4:0] id; logic user; logic [31:0] addr; logic [7:0] length; logic [2:0] size; logic [1:0] burst; logic lock; logic [3:0] cache; logic [2:0] prot; logic [3:0] qos; logic [3:0] region; }
    _Cache_inst0_nasti_ar_data;
  wire _Cache_inst0_nasti_r_ready;
  wire _MemArbiter_inst0_icache_aw_ready;
  wire _MemArbiter_inst0_icache_w_ready;
  wire _MemArbiter_inst0_icache_b_valid;
  wire struct packed {logic [1:0] resp; logic [4:0] id; logic user; }
    _MemArbiter_inst0_icache_b_data;
  wire _MemArbiter_inst0_icache_ar_ready;
  wire _MemArbiter_inst0_icache_r_valid;
  wire
    struct packed {logic [1:0] resp; logic [4:0] id; logic user; logic [63:0] data; logic last; }
    _MemArbiter_inst0_icache_r_data;
  wire _MemArbiter_inst0_dcache_aw_ready;
  wire _MemArbiter_inst0_dcache_w_ready;
  wire _MemArbiter_inst0_dcache_b_valid;
  wire struct packed {logic [1:0] resp; logic [4:0] id; logic user; }
    _MemArbiter_inst0_dcache_b_data;
  wire _MemArbiter_inst0_dcache_ar_ready;
  wire _MemArbiter_inst0_dcache_r_valid;
  wire
    struct packed {logic [1:0] resp; logic [4:0] id; logic user; logic [63:0] data; logic last; }
    _MemArbiter_inst0_dcache_r_data;
  wire struct packed {logic valid; struct packed {logic [31:0] data; } data; }
    _Cache_inst1_cpu_resp;
  wire _Cache_inst1_nasti_aw_valid;
  wire
    struct packed {logic [4:0] id; logic user; logic [31:0] addr; logic [7:0] length; logic [2:0] size; logic [1:0] burst; logic lock; logic [3:0] cache; logic [2:0] prot; logic [3:0] qos; logic [3:0] region; }
    _Cache_inst1_nasti_aw_data;
  wire _Cache_inst1_nasti_w_valid;
  wire
    struct packed {logic [4:0] id; logic [7:0] strb; logic user; logic [63:0] data; logic last; }
    _Cache_inst1_nasti_w_data;
  wire _Cache_inst1_nasti_b_ready;
  wire _Cache_inst1_nasti_ar_valid;
  wire
    struct packed {logic [4:0] id; logic user; logic [31:0] addr; logic [7:0] length; logic [2:0] size; logic [1:0] burst; logic lock; logic [3:0] cache; logic [2:0] prot; logic [3:0] qos; logic [3:0] region; }
    _Cache_inst1_nasti_ar_data;
  wire _Cache_inst1_nasti_r_ready;
  Cache Cache_inst1 (
    .cpu_abort      (_Core_inst0_dcache_abort),
    .cpu_req        (_Core_inst0_dcache_req),
    .nasti_aw_ready (_MemArbiter_inst0_dcache_aw_ready),
    .nasti_w_ready  (_MemArbiter_inst0_dcache_w_ready),
    .nasti_b_valid  (_MemArbiter_inst0_dcache_b_valid),
    .nasti_b_data   (_MemArbiter_inst0_dcache_b_data),
    .nasti_ar_ready (_MemArbiter_inst0_dcache_ar_ready),
    .nasti_r_valid  (_MemArbiter_inst0_dcache_r_valid),
    .nasti_r_data   (_MemArbiter_inst0_dcache_r_data),
    .CLK            (CLK),
    .RESET          (RESET),
    .cpu_resp       (_Cache_inst1_cpu_resp),
    .nasti_aw_valid (_Cache_inst1_nasti_aw_valid),
    .nasti_aw_data  (_Cache_inst1_nasti_aw_data),
    .nasti_w_valid  (_Cache_inst1_nasti_w_valid),
    .nasti_w_data   (_Cache_inst1_nasti_w_data),
    .nasti_b_ready  (_Cache_inst1_nasti_b_ready),
    .nasti_ar_valid (_Cache_inst1_nasti_ar_valid),
    .nasti_ar_data  (_Cache_inst1_nasti_ar_data),
    .nasti_r_ready  (_Cache_inst1_nasti_r_ready)
  );
  MemArbiter MemArbiter_inst0 (
    .icache_aw_valid (_Cache_inst0_nasti_aw_valid),
    .icache_aw_data  (_Cache_inst0_nasti_aw_data),
    .icache_w_valid  (_Cache_inst0_nasti_w_valid),
    .icache_w_data   (_Cache_inst0_nasti_w_data),
    .icache_b_ready  (_Cache_inst0_nasti_b_ready),
    .icache_ar_valid (_Cache_inst0_nasti_ar_valid),
    .icache_ar_data  (_Cache_inst0_nasti_ar_data),
    .icache_r_ready  (_Cache_inst0_nasti_r_ready),
    .dcache_aw_valid (_Cache_inst1_nasti_aw_valid),
    .dcache_aw_data  (_Cache_inst1_nasti_aw_data),
    .dcache_w_valid  (_Cache_inst1_nasti_w_valid),
    .dcache_w_data   (_Cache_inst1_nasti_w_data),
    .dcache_b_ready  (_Cache_inst1_nasti_b_ready),
    .dcache_ar_valid (_Cache_inst1_nasti_ar_valid),
    .dcache_ar_data  (_Cache_inst1_nasti_ar_data),
    .dcache_r_ready  (_Cache_inst1_nasti_r_ready),
    .nasti_aw_ready  (nasti_aw_ready),
    .nasti_w_ready   (nasti_w_ready),
    .nasti_b_valid   (nasti_b_valid),
    .nasti_b_data    (nasti_b_data),
    .nasti_ar_ready  (nasti_ar_ready),
    .nasti_r_valid   (nasti_r_valid),
    .nasti_r_data    (nasti_r_data),
    .CLK             (CLK),
    .RESET           (RESET),
    .icache_aw_ready (_MemArbiter_inst0_icache_aw_ready),
    .icache_w_ready  (_MemArbiter_inst0_icache_w_ready),
    .icache_b_valid  (_MemArbiter_inst0_icache_b_valid),
    .icache_b_data   (_MemArbiter_inst0_icache_b_data),
    .icache_ar_ready (_MemArbiter_inst0_icache_ar_ready),
    .icache_r_valid  (_MemArbiter_inst0_icache_r_valid),
    .icache_r_data   (_MemArbiter_inst0_icache_r_data),
    .dcache_aw_ready (_MemArbiter_inst0_dcache_aw_ready),
    .dcache_w_ready  (_MemArbiter_inst0_dcache_w_ready),
    .dcache_b_valid  (_MemArbiter_inst0_dcache_b_valid),
    .dcache_b_data   (_MemArbiter_inst0_dcache_b_data),
    .dcache_ar_ready (_MemArbiter_inst0_dcache_ar_ready),
    .dcache_r_valid  (_MemArbiter_inst0_dcache_r_valid),
    .dcache_r_data   (_MemArbiter_inst0_dcache_r_data),
    .nasti_aw_valid  (nasti_aw_valid),
    .nasti_aw_data   (nasti_aw_data),
    .nasti_w_valid   (nasti_w_valid),
    .nasti_w_data    (nasti_w_data),
    .nasti_b_ready   (nasti_b_ready),
    .nasti_ar_valid  (nasti_ar_valid),
    .nasti_ar_data   (nasti_ar_data),
    .nasti_r_ready   (nasti_r_ready)
  );
  Cache Cache_inst0 (
    .cpu_abort      (_Core_inst0_icache_abort),
    .cpu_req        (_Core_inst0_icache_req),
    .nasti_aw_ready (_MemArbiter_inst0_icache_aw_ready),
    .nasti_w_ready  (_MemArbiter_inst0_icache_w_ready),
    .nasti_b_valid  (_MemArbiter_inst0_icache_b_valid),
    .nasti_b_data   (_MemArbiter_inst0_icache_b_data),
    .nasti_ar_ready (_MemArbiter_inst0_icache_ar_ready),
    .nasti_r_valid  (_MemArbiter_inst0_icache_r_valid),
    .nasti_r_data   (_MemArbiter_inst0_icache_r_data),
    .CLK            (CLK),
    .RESET          (RESET),
    .cpu_resp       (_Cache_inst0_cpu_resp),
    .nasti_aw_valid (_Cache_inst0_nasti_aw_valid),
    .nasti_aw_data  (_Cache_inst0_nasti_aw_data),
    .nasti_w_valid  (_Cache_inst0_nasti_w_valid),
    .nasti_w_data   (_Cache_inst0_nasti_w_data),
    .nasti_b_ready  (_Cache_inst0_nasti_b_ready),
    .nasti_ar_valid (_Cache_inst0_nasti_ar_valid),
    .nasti_ar_data  (_Cache_inst0_nasti_ar_data),
    .nasti_r_ready  (_Cache_inst0_nasti_r_ready)
  );
  Core Core_inst0 (
    .host_fromhost (host_fromhost),
    .icache_resp   (_Cache_inst0_cpu_resp),
    .dcache_resp   (_Cache_inst1_cpu_resp),
    .CLK           (CLK),
    .RESET         (RESET),
    .host_tohost   (host_tohost),
    .icache_abort  (_Core_inst0_icache_abort),
    .icache_req    (_Core_inst0_icache_req),
    .dcache_abort  (_Core_inst0_dcache_abort),
    .dcache_req    (_Core_inst0_dcache_req)
  );
endmodule

