module simple_wrap_cast(
  input  I,
  output O);

  assign O = I;	// <stdin>:3:5
endmodule

