module coreir_term #(
    parameter width = 1
) (
    input [width-1:0] in
);

endmodule

module MonitorWrapper (
    input [7:0] arr_0,
    input [7:0] arr_1,
    input [7:0] arr_10,
    input [7:0] arr_11,
    input [7:0] arr_12,
    input [7:0] arr_13,
    input [7:0] arr_14,
    input [7:0] arr_15,
    input [7:0] arr_16,
    input [7:0] arr_17,
    input [7:0] arr_18,
    input [7:0] arr_19,
    input [7:0] arr_2,
    input [7:0] arr_20,
    input [7:0] arr_21,
    input [7:0] arr_22,
    input [7:0] arr_23,
    input [7:0] arr_24,
    input [7:0] arr_25,
    input [7:0] arr_26,
    input [7:0] arr_27,
    input [7:0] arr_28,
    input [7:0] arr_29,
    input [7:0] arr_3,
    input [7:0] arr_30,
    input [7:0] arr_31,
    input [7:0] arr_32,
    input [7:0] arr_33,
    input [7:0] arr_34,
    input [7:0] arr_35,
    input [7:0] arr_36,
    input [7:0] arr_37,
    input [7:0] arr_38,
    input [7:0] arr_39,
    input [7:0] arr_4,
    input [7:0] arr_40,
    input [7:0] arr_41,
    input [7:0] arr_42,
    input [7:0] arr_43,
    input [7:0] arr_44,
    input [7:0] arr_45,
    input [7:0] arr_46,
    input [7:0] arr_47,
    input [7:0] arr_48,
    input [7:0] arr_49,
    input [7:0] arr_5,
    input [7:0] arr_50,
    input [7:0] arr_51,
    input [7:0] arr_52,
    input [7:0] arr_53,
    input [7:0] arr_54,
    input [7:0] arr_55,
    input [7:0] arr_56,
    input [7:0] arr_57,
    input [7:0] arr_58,
    input [7:0] arr_59,
    input [7:0] arr_6,
    input [7:0] arr_60,
    input [7:0] arr_61,
    input [7:0] arr_62,
    input [7:0] arr_63,
    input [7:0] arr_7,
    input [7:0] arr_8,
    input [7:0] arr_9
);
coreir_term #(
    .width(8)
) term_inst0 (
    .in(arr_0)
);
coreir_term #(
    .width(8)
) term_inst1 (
    .in(arr_1)
);
coreir_term #(
    .width(8)
) term_inst10 (
    .in(arr_10)
);
coreir_term #(
    .width(8)
) term_inst11 (
    .in(arr_11)
);
coreir_term #(
    .width(8)
) term_inst12 (
    .in(arr_12)
);
coreir_term #(
    .width(8)
) term_inst13 (
    .in(arr_13)
);
coreir_term #(
    .width(8)
) term_inst14 (
    .in(arr_14)
);
coreir_term #(
    .width(8)
) term_inst15 (
    .in(arr_15)
);
coreir_term #(
    .width(8)
) term_inst16 (
    .in(arr_16)
);
coreir_term #(
    .width(8)
) term_inst17 (
    .in(arr_17)
);
coreir_term #(
    .width(8)
) term_inst18 (
    .in(arr_18)
);
coreir_term #(
    .width(8)
) term_inst19 (
    .in(arr_19)
);
coreir_term #(
    .width(8)
) term_inst2 (
    .in(arr_2)
);
coreir_term #(
    .width(8)
) term_inst20 (
    .in(arr_20)
);
coreir_term #(
    .width(8)
) term_inst21 (
    .in(arr_21)
);
coreir_term #(
    .width(8)
) term_inst22 (
    .in(arr_22)
);
coreir_term #(
    .width(8)
) term_inst23 (
    .in(arr_23)
);
coreir_term #(
    .width(8)
) term_inst24 (
    .in(arr_24)
);
coreir_term #(
    .width(8)
) term_inst25 (
    .in(arr_25)
);
coreir_term #(
    .width(8)
) term_inst26 (
    .in(arr_26)
);
coreir_term #(
    .width(8)
) term_inst27 (
    .in(arr_27)
);
coreir_term #(
    .width(8)
) term_inst28 (
    .in(arr_28)
);
coreir_term #(
    .width(8)
) term_inst29 (
    .in(arr_29)
);
coreir_term #(
    .width(8)
) term_inst3 (
    .in(arr_3)
);
coreir_term #(
    .width(8)
) term_inst30 (
    .in(arr_30)
);
coreir_term #(
    .width(8)
) term_inst31 (
    .in(arr_31)
);
coreir_term #(
    .width(8)
) term_inst32 (
    .in(arr_32)
);
coreir_term #(
    .width(8)
) term_inst33 (
    .in(arr_33)
);
coreir_term #(
    .width(8)
) term_inst34 (
    .in(arr_34)
);
coreir_term #(
    .width(8)
) term_inst35 (
    .in(arr_35)
);
coreir_term #(
    .width(8)
) term_inst36 (
    .in(arr_36)
);
coreir_term #(
    .width(8)
) term_inst37 (
    .in(arr_37)
);
coreir_term #(
    .width(8)
) term_inst38 (
    .in(arr_38)
);
coreir_term #(
    .width(8)
) term_inst39 (
    .in(arr_39)
);
coreir_term #(
    .width(8)
) term_inst4 (
    .in(arr_4)
);
coreir_term #(
    .width(8)
) term_inst40 (
    .in(arr_40)
);
coreir_term #(
    .width(8)
) term_inst41 (
    .in(arr_41)
);
coreir_term #(
    .width(8)
) term_inst42 (
    .in(arr_42)
);
coreir_term #(
    .width(8)
) term_inst43 (
    .in(arr_43)
);
coreir_term #(
    .width(8)
) term_inst44 (
    .in(arr_44)
);
coreir_term #(
    .width(8)
) term_inst45 (
    .in(arr_45)
);
coreir_term #(
    .width(8)
) term_inst46 (
    .in(arr_46)
);
coreir_term #(
    .width(8)
) term_inst47 (
    .in(arr_47)
);
coreir_term #(
    .width(8)
) term_inst48 (
    .in(arr_48)
);
coreir_term #(
    .width(8)
) term_inst49 (
    .in(arr_49)
);
coreir_term #(
    .width(8)
) term_inst5 (
    .in(arr_5)
);
coreir_term #(
    .width(8)
) term_inst50 (
    .in(arr_50)
);
coreir_term #(
    .width(8)
) term_inst51 (
    .in(arr_51)
);
coreir_term #(
    .width(8)
) term_inst52 (
    .in(arr_52)
);
coreir_term #(
    .width(8)
) term_inst53 (
    .in(arr_53)
);
coreir_term #(
    .width(8)
) term_inst54 (
    .in(arr_54)
);
coreir_term #(
    .width(8)
) term_inst55 (
    .in(arr_55)
);
coreir_term #(
    .width(8)
) term_inst56 (
    .in(arr_56)
);
coreir_term #(
    .width(8)
) term_inst57 (
    .in(arr_57)
);
coreir_term #(
    .width(8)
) term_inst58 (
    .in(arr_58)
);
coreir_term #(
    .width(8)
) term_inst59 (
    .in(arr_59)
);
coreir_term #(
    .width(8)
) term_inst6 (
    .in(arr_6)
);
coreir_term #(
    .width(8)
) term_inst60 (
    .in(arr_60)
);
coreir_term #(
    .width(8)
) term_inst61 (
    .in(arr_61)
);
coreir_term #(
    .width(8)
) term_inst62 (
    .in(arr_62)
);
coreir_term #(
    .width(8)
) term_inst63 (
    .in(arr_63)
);
coreir_term #(
    .width(8)
) term_inst7 (
    .in(arr_7)
);
coreir_term #(
    .width(8)
) term_inst8 (
    .in(arr_8)
);
coreir_term #(
    .width(8)
) term_inst9 (
    .in(arr_9)
);

monitor #(.WIDTH(8), .DEPTH(64)) monitor_inst(.arr('{arr_63, arr_62, arr_61, arr_60, arr_59, arr_58, arr_57, arr_56, arr_55, arr_54, arr_53, arr_52, arr_51, arr_50, arr_49, arr_48, arr_47, arr_46, arr_45, arr_44, arr_43, arr_42, arr_41, arr_40, arr_39, arr_38, arr_37, arr_36, arr_35, arr_34, arr_33, arr_32, arr_31, arr_30, arr_29, arr_28, arr_27, arr_26, arr_25, arr_24, arr_23, arr_22, arr_21, arr_20, arr_19, arr_18, arr_17, arr_16, arr_15, arr_14, arr_13, arr_12, arr_11, arr_10, arr_9, arr_8, arr_7, arr_6, arr_5, arr_4, arr_3, arr_2, arr_1, arr_0}));
                    
endmodule

