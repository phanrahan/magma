module feedthrough(
  input  I,
  output O);

  assign O = I;	// <stdin>:3:5
endmodule

