module simple_aggregates_array(
  input  [7:0][15:0] a,
  output [7:0][15:0] y);

  assign y = {{a[3'h3]}, {a[3'h2]}, {a[3'h1]}, {a[3'h0]}, {a[3'h7]}, {a[3'h6]}, {a[3'h5]}, {a[3'h4]}};	// <stdin>:3:14, :4:14, :5:14, :6:14, :7:15, :8:15, :9:15, :10:15, :11:10, :12:10, :13:10, :14:10, :15:10, :16:10, :17:10, :18:10, :19:10, :20:5
endmodule

