// external module simple_verilog_defn

module simple_verilog_defn_wrapper(	// <stdin>:2:1
  input  I,
  output O);

  simple_verilog_defn simple_verilog_defn_inst0 (	// <stdin>:3:10
    .I (I),
    .O (O)
  );
endmodule

