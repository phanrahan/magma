// external module simple_decl

module simple_decl_external(	// <stdin>:2:1
  input  I,
  output O);

  simple_decl simple_decl_inst0 (	// <stdin>:3:10
    .I (I),
    .O (O)
  );
endmodule

