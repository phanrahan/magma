module feedthrough(	// <stdin>:1:1
  input  I,
  output O);

  assign O = I;	// <stdin>:2:5
endmodule

