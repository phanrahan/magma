module main (output [1:0] LED, input [1:0] SWITCH);
assign LED = SWITCH;
endmodule

