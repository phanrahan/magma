module mod0 #(parameter KRATOS_INSTANCE_ID = 32'hDEADBEEF)
(
    input I
);

endmodule   // mod
