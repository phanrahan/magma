module Mux6xTuplex_Bits8_y_Bit(
  input  struct packed {logic [7:0] x; logic y; } I0, I1, I2, I3, I4, I5,
  input  [2:0]                                    S,
  output struct packed {logic [7:0] x; logic y; } O);

  wire [7:0] _T = I0.x;	// <stdin>:3:10
  wire [7:0] _T_0 = I0.x;	// <stdin>:5:10
  wire [7:0] _T_1 = I0.x;	// <stdin>:7:10
  wire [7:0] _T_2 = I0.x;	// <stdin>:9:10
  wire [7:0] _T_3 = I0.x;	// <stdin>:11:10
  wire [7:0] _T_4 = I0.x;	// <stdin>:13:11
  wire [7:0] _T_5 = I0.x;	// <stdin>:15:11
  wire [7:0] _T_6 = I0.x;	// <stdin>:17:11
  wire [7:0] _T_7 = I1.x;	// <stdin>:21:11
  wire [7:0] _T_8 = I1.x;	// <stdin>:23:11
  wire [7:0] _T_9 = I1.x;	// <stdin>:25:11
  wire [7:0] _T_10 = I1.x;	// <stdin>:27:11
  wire [7:0] _T_11 = I1.x;	// <stdin>:29:11
  wire [7:0] _T_12 = I1.x;	// <stdin>:31:11
  wire [7:0] _T_13 = I1.x;	// <stdin>:33:11
  wire [7:0] _T_14 = I1.x;	// <stdin>:35:11
  wire [7:0] _T_15 = I2.x;	// <stdin>:39:11
  wire [7:0] _T_16 = I2.x;	// <stdin>:41:11
  wire [7:0] _T_17 = I2.x;	// <stdin>:43:11
  wire [7:0] _T_18 = I2.x;	// <stdin>:45:11
  wire [7:0] _T_19 = I2.x;	// <stdin>:47:11
  wire [7:0] _T_20 = I2.x;	// <stdin>:49:11
  wire [7:0] _T_21 = I2.x;	// <stdin>:51:11
  wire [7:0] _T_22 = I2.x;	// <stdin>:53:11
  wire [7:0] _T_23 = I3.x;	// <stdin>:57:11
  wire [7:0] _T_24 = I3.x;	// <stdin>:59:11
  wire [7:0] _T_25 = I3.x;	// <stdin>:61:11
  wire [7:0] _T_26 = I3.x;	// <stdin>:63:11
  wire [7:0] _T_27 = I3.x;	// <stdin>:65:11
  wire [7:0] _T_28 = I3.x;	// <stdin>:67:11
  wire [7:0] _T_29 = I3.x;	// <stdin>:69:11
  wire [7:0] _T_30 = I3.x;	// <stdin>:71:11
  wire [7:0] _T_31 = I4.x;	// <stdin>:75:11
  wire [7:0] _T_32 = I4.x;	// <stdin>:77:11
  wire [7:0] _T_33 = I4.x;	// <stdin>:79:11
  wire [7:0] _T_34 = I4.x;	// <stdin>:81:11
  wire [7:0] _T_35 = I4.x;	// <stdin>:83:11
  wire [7:0] _T_36 = I4.x;	// <stdin>:85:11
  wire [7:0] _T_37 = I4.x;	// <stdin>:87:11
  wire [7:0] _T_38 = I4.x;	// <stdin>:89:11
  wire [7:0] _T_39 = I5.x;	// <stdin>:93:11
  wire [7:0] _T_40 = I5.x;	// <stdin>:95:11
  wire [7:0] _T_41 = I5.x;	// <stdin>:97:11
  wire [7:0] _T_42 = I5.x;	// <stdin>:99:11
  wire [7:0] _T_43 = I5.x;	// <stdin>:101:11
  wire [7:0] _T_44 = I5.x;	// <stdin>:103:12
  wire [7:0] _T_45 = I5.x;	// <stdin>:105:12
  wire [7:0] _T_46 = I5.x;	// <stdin>:107:12
  wire [8:0] _tmp = {I5.y, _T_46[7], _T_45[6], _T_44[5], _T_43[4], _T_42[3], _T_41[2], _T_40[1], _T_39[0]};	// <stdin>:94:11, :96:11, :98:11, :100:11, :102:11, :104:12, :106:12, :108:12, :109:12, :110:12
  wire [8:0] _tmp_50 = {I4.y, _T_38[7], _T_37[6], _T_36[5], _T_35[4], _T_34[3], _T_33[2], _T_32[1], _T_31[0]};	// <stdin>:76:11, :78:11, :80:11, :82:11, :84:11, :86:11, :88:11, :90:11, :91:11, :92:11
  wire [8:0] _tmp_51 = {I3.y, _T_30[7], _T_29[6], _T_28[5], _T_27[4], _T_26[3], _T_25[2], _T_24[1], _T_23[0]};	// <stdin>:58:11, :60:11, :62:11, :64:11, :66:11, :68:11, :70:11, :72:11, :73:11, :74:11
  wire [8:0] _tmp_52 = {I2.y, _T_22[7], _T_21[6], _T_20[5], _T_19[4], _T_18[3], _T_17[2], _T_16[1], _T_15[0]};	// <stdin>:40:11, :42:11, :44:11, :46:11, :48:11, :50:11, :52:11, :54:11, :55:11, :56:11
  wire [8:0] _tmp_53 = {I1.y, _T_14[7], _T_13[6], _T_12[5], _T_11[4], _T_10[3], _T_9[2], _T_8[1], _T_7[0]};	// <stdin>:22:11, :24:11, :26:11, :28:11, :30:11, :32:11, :34:11, :36:11, :37:11, :38:11
  wire [8:0] _tmp_54 = {I0.y, _T_6[7], _T_5[6], _T_4[5], _T_3[4], _T_2[3], _T_1[2], _T_0[1], _T[0]};	// <stdin>:4:10, :6:10, :8:10, :10:10, :12:10, :14:11, :16:11, :18:11, :19:11, :20:11
  wire [5:0][8:0] _tmp_55 = {{_tmp}, {_tmp_50}, {_tmp_51}, {_tmp_52}, {_tmp_53}, {_tmp_54}};	// <stdin>:111:12
  wire struct packed {logic [5:0][8:0] data; logic [2:0] sel; } _T_47 = '{data: _tmp_55, sel: S};	// <stdin>:4:10, :6:10, :8:10, :10:10, :12:10, :14:11, :16:11, :18:11, :19:11, :22:11, :24:11, :26:11, :28:11, :30:11, :32:11, :34:11, :36:11, :37:11, :40:11, :42:11, :44:11, :46:11, :48:11, :50:11, :52:11, :54:11, :55:11, :58:11, :60:11, :62:11, :64:11, :66:11, :68:11, :70:11, :72:11, :73:11, :76:11, :78:11, :80:11, :82:11, :84:11, :86:11, :88:11, :90:11, :91:11, :94:11, :96:11, :98:11, :100:11, :102:11, :104:12, :106:12, :108:12, :109:12, :112:12
  wire [8:0] _T_48 = _T_47.data[_T_47.sel];	// <stdin>:113:12, :114:12, :115:12
  wire struct packed {logic [7:0] x; logic y; } _T_49 = '{x: (_T_48[7:0]), y: (_T_48[8])};	// <stdin>:116:12, :117:12, :118:12
  assign O = _T_49;	// <stdin>:119:5
endmodule

