module simple_inline_verilog(	// <stdin>:1:1
  input  I,
  output O);

  
  	// This is 'a' "comment".	// <stdin>:3:5
  assign O = I;	// <stdin>:4:5
endmodule

