module return_magma_named_tuple (input [1:0] I, output  O_x, output  O_y);
assign O_x = I[0];
assign O_y = I[1];
endmodule

