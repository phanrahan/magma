module main (output [7:0] LED, input [7:0] SWITCH);
assign LED = SWITCH;
endmodule

