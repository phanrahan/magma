module simple_inline_verilog(
  input  I,
  output O
);


  	// This is 'a' "comment".
  assign O = I;
endmodule

