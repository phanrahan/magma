module main (input  I, output  O);
assign O = I;
endmodule

