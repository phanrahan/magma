// Module `PRWDWUWSWCDGH_V` defined externally
module corebit_const #(
    parameter value = 1
) (
    output out
);
  assign out = value;
endmodule

module Top (
    inout pad
);
wire PRWDWUWSWCDGH_V_inst0_C;
wire PRWDWUWSWCDGH_V_inst0_DS0;
wire PRWDWUWSWCDGH_V_inst0_DS1;
wire PRWDWUWSWCDGH_V_inst0_DS2;
wire PRWDWUWSWCDGH_V_inst0_I;
wire PRWDWUWSWCDGH_V_inst0_IE;
wire PRWDWUWSWCDGH_V_inst0_OEN;
wire PRWDWUWSWCDGH_V_inst0_PAD;
wire PRWDWUWSWCDGH_V_inst0_PU;
wire PRWDWUWSWCDGH_V_inst0_PD;
wire PRWDWUWSWCDGH_V_inst0_ST;
wire PRWDWUWSWCDGH_V_inst0_SL;
wire PRWDWUWSWCDGH_V_inst0_RTE;
wire bit_const_0_None_out;
assign PRWDWUWSWCDGH_V_inst0_DS0 = bit_const_0_None_out;
assign PRWDWUWSWCDGH_V_inst0_DS1 = bit_const_0_None_out;
assign PRWDWUWSWCDGH_V_inst0_DS2 = bit_const_0_None_out;
assign PRWDWUWSWCDGH_V_inst0_I = bit_const_0_None_out;
assign PRWDWUWSWCDGH_V_inst0_IE = bit_const_0_None_out;
assign PRWDWUWSWCDGH_V_inst0_OEN = bit_const_0_None_out;
assign PRWDWUWSWCDGH_V_inst0_PU = bit_const_0_None_out;
assign PRWDWUWSWCDGH_V_inst0_PD = bit_const_0_None_out;
assign PRWDWUWSWCDGH_V_inst0_ST = bit_const_0_None_out;
assign PRWDWUWSWCDGH_V_inst0_SL = bit_const_0_None_out;
assign PRWDWUWSWCDGH_V_inst0_RTE = bit_const_0_None_out;
PRWDWUWSWCDGH_V PRWDWUWSWCDGH_V_inst0 (
    .C(PRWDWUWSWCDGH_V_inst0_C),
    .DS0(PRWDWUWSWCDGH_V_inst0_DS0),
    .DS1(PRWDWUWSWCDGH_V_inst0_DS1),
    .DS2(PRWDWUWSWCDGH_V_inst0_DS2),
    .I(PRWDWUWSWCDGH_V_inst0_I),
    .IE(PRWDWUWSWCDGH_V_inst0_IE),
    .OEN(PRWDWUWSWCDGH_V_inst0_OEN),
    .PAD(PRWDWUWSWCDGH_V_inst0_PAD),
    .PU(PRWDWUWSWCDGH_V_inst0_PU),
    .PD(PRWDWUWSWCDGH_V_inst0_PD),
    .ST(PRWDWUWSWCDGH_V_inst0_ST),
    .SL(PRWDWUWSWCDGH_V_inst0_SL),
    .RTE(PRWDWUWSWCDGH_V_inst0_RTE)
);
corebit_const #(
    .value(1'b0)
) bit_const_0_None (
    .out(bit_const_0_None_out)
);
assign PRWDWUWSWCDGH_V_inst0_PAD = pad;
endmodule

