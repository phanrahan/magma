module mod1 #(parameter KRATOS_INSTANCE_ID = 'h1)
(
    input I
);

endmodule   // mod
