module file(
  input                                                        CLK, ASYNCRESET,
  input  [7:0]                                                 file_read_0_addr,
  input  [7:0]                                                 file_read_1_addr,
  input  struct packed {logic [31:0] data; logic [7:0] addr; } write_0,
  input                                                        write_0_en,
  output [31:0]                                                file_read_0_data,
  output [31:0]                                                file_read_1_data);

  wire [31:0] _T;	// <stdin>:3081:13
  wire [31:0] _T_0;	// <stdin>:2298:13
  wire [31:0] _T_1;	// <stdin>:2290:13
  wire [31:0] _T_2;	// <stdin>:2282:13
  wire [31:0] _T_3;	// <stdin>:2274:13
  wire [31:0] _T_4;	// <stdin>:2266:13
  wire [31:0] _T_5;	// <stdin>:2258:13
  wire [31:0] _T_6;	// <stdin>:2250:13
  wire [31:0] _T_7;	// <stdin>:2242:13
  wire [31:0] _T_8;	// <stdin>:2234:13
  wire [31:0] _T_9;	// <stdin>:2226:13
  wire [31:0] _T_10;	// <stdin>:2218:13
  wire [31:0] _T_11;	// <stdin>:2210:13
  wire [31:0] _T_12;	// <stdin>:2202:13
  wire [31:0] _T_13;	// <stdin>:2194:13
  wire [31:0] _T_14;	// <stdin>:2186:13
  wire [31:0] _T_15;	// <stdin>:2178:13
  wire [31:0] _T_16;	// <stdin>:2170:13
  wire [31:0] _T_17;	// <stdin>:2162:13
  wire [31:0] _T_18;	// <stdin>:2154:13
  wire [31:0] _T_19;	// <stdin>:2146:13
  wire [31:0] _T_20;	// <stdin>:2138:13
  wire [31:0] _T_21;	// <stdin>:2130:13
  wire [31:0] _T_22;	// <stdin>:2122:13
  wire [31:0] _T_23;	// <stdin>:2114:13
  wire [31:0] _T_24;	// <stdin>:2106:13
  wire [31:0] _T_25;	// <stdin>:2098:13
  wire [31:0] _T_26;	// <stdin>:2090:13
  wire [31:0] _T_27;	// <stdin>:2082:13
  wire [31:0] _T_28;	// <stdin>:2074:13
  wire [31:0] _T_29;	// <stdin>:2066:13
  wire [31:0] _T_30;	// <stdin>:2058:13
  wire [31:0] _T_31;	// <stdin>:2050:13
  wire [31:0] _T_32;	// <stdin>:2042:13
  wire [31:0] _T_33;	// <stdin>:2034:13
  wire [31:0] _T_34;	// <stdin>:2026:13
  wire [31:0] _T_35;	// <stdin>:2018:13
  wire [31:0] _T_36;	// <stdin>:2010:13
  wire [31:0] _T_37;	// <stdin>:2002:13
  wire [31:0] _T_38;	// <stdin>:1994:13
  wire [31:0] _T_39;	// <stdin>:1986:13
  wire [31:0] _T_40;	// <stdin>:1978:13
  wire [31:0] _T_41;	// <stdin>:1970:13
  wire [31:0] _T_42;	// <stdin>:1962:13
  wire [31:0] _T_43;	// <stdin>:1954:13
  wire [31:0] _T_44;	// <stdin>:1946:13
  wire [31:0] _T_45;	// <stdin>:1938:13
  wire [31:0] _T_46;	// <stdin>:1930:13
  wire [31:0] _T_47;	// <stdin>:1922:13
  wire [31:0] _T_48;	// <stdin>:1914:13
  wire [31:0] _T_49;	// <stdin>:1906:13
  wire [31:0] _T_50;	// <stdin>:1898:13
  wire [31:0] _T_51;	// <stdin>:1890:13
  wire [31:0] _T_52;	// <stdin>:1882:13
  wire [31:0] _T_53;	// <stdin>:1874:13
  wire [31:0] _T_54;	// <stdin>:1866:13
  wire [31:0] _T_55;	// <stdin>:1858:13
  wire [31:0] _T_56;	// <stdin>:1850:13
  wire [31:0] _T_57;	// <stdin>:1842:13
  wire [31:0] _T_58;	// <stdin>:1834:13
  wire [31:0] _T_59;	// <stdin>:1826:13
  wire [31:0] _T_60;	// <stdin>:1818:13
  wire [31:0] _T_61;	// <stdin>:1810:13
  wire [31:0] _T_62;	// <stdin>:1802:13
  wire [31:0] _T_63;	// <stdin>:1794:13
  wire [31:0] _T_64;	// <stdin>:1786:13
  wire [31:0] _T_65;	// <stdin>:1778:13
  wire [31:0] _T_66;	// <stdin>:1770:13
  wire [31:0] _T_67;	// <stdin>:1762:13
  wire [31:0] _T_68;	// <stdin>:1754:13
  wire [31:0] _T_69;	// <stdin>:1746:13
  wire [31:0] _T_70;	// <stdin>:1738:13
  wire [31:0] _T_71;	// <stdin>:1730:13
  wire [31:0] _T_72;	// <stdin>:1722:13
  wire [31:0] _T_73;	// <stdin>:1714:13
  wire [31:0] _T_74;	// <stdin>:1706:13
  wire [31:0] _T_75;	// <stdin>:1698:13
  wire [31:0] _T_76;	// <stdin>:1690:13
  wire [31:0] _T_77;	// <stdin>:1682:13
  wire [31:0] _T_78;	// <stdin>:1674:13
  wire [31:0] _T_79;	// <stdin>:1666:13
  wire [31:0] _T_80;	// <stdin>:1658:13
  wire [31:0] _T_81;	// <stdin>:1650:13
  wire [31:0] _T_82;	// <stdin>:1642:13
  wire [31:0] _T_83;	// <stdin>:1634:13
  wire [31:0] _T_84;	// <stdin>:1626:13
  wire [31:0] _T_85;	// <stdin>:1618:13
  wire [31:0] _T_86;	// <stdin>:1610:13
  wire [31:0] _T_87;	// <stdin>:1602:13
  wire [31:0] _T_88;	// <stdin>:1594:13
  wire [31:0] _T_89;	// <stdin>:1586:13
  wire [31:0] _T_90;	// <stdin>:1578:13
  wire [31:0] _T_91;	// <stdin>:1570:13
  wire [31:0] _T_92;	// <stdin>:1562:13
  wire [31:0] _T_93;	// <stdin>:1554:13
  wire [31:0] _T_94;	// <stdin>:1546:13
  wire [31:0] _T_95;	// <stdin>:1538:13
  wire [31:0] _T_96;	// <stdin>:1530:13
  wire [31:0] _T_97;	// <stdin>:1522:13
  wire [31:0] _T_98;	// <stdin>:1514:13
  wire [31:0] _T_99;	// <stdin>:1506:13
  wire [31:0] _T_100;	// <stdin>:1498:13
  wire [31:0] _T_101;	// <stdin>:1490:13
  wire [31:0] _T_102;	// <stdin>:1482:13
  wire [31:0] _T_103;	// <stdin>:1474:13
  wire [31:0] _T_104;	// <stdin>:1466:13
  wire [31:0] _T_105;	// <stdin>:1458:13
  wire [31:0] _T_106;	// <stdin>:1450:13
  wire [31:0] _T_107;	// <stdin>:1442:13
  wire [31:0] _T_108;	// <stdin>:1434:13
  wire [31:0] _T_109;	// <stdin>:1426:13
  wire [31:0] _T_110;	// <stdin>:1418:13
  wire [31:0] _T_111;	// <stdin>:1410:13
  wire [31:0] _T_112;	// <stdin>:1402:13
  wire [31:0] _T_113;	// <stdin>:1394:12
  wire [31:0] _T_114;	// <stdin>:1386:12
  wire [31:0] _T_115;	// <stdin>:1378:12
  wire [31:0] _T_116;	// <stdin>:1370:12
  wire [31:0] _T_117;	// <stdin>:1362:12
  wire [31:0] _T_118;	// <stdin>:1354:12
  wire [31:0] _T_119;	// <stdin>:1346:12
  wire [31:0] _T_120;	// <stdin>:1338:12
  wire [31:0] _T_121;	// <stdin>:1330:12
  wire [31:0] _T_122;	// <stdin>:1322:12
  wire [31:0] _T_123;	// <stdin>:1314:12
  wire [31:0] _T_124;	// <stdin>:1306:12
  wire [31:0] _T_125;	// <stdin>:1298:12
  wire [31:0] _T_126;	// <stdin>:1290:12
  wire [31:0] _T_127;	// <stdin>:1282:12
  wire [31:0] _T_128;	// <stdin>:1274:12
  wire [31:0] _T_129;	// <stdin>:1266:12
  wire [31:0] _T_130;	// <stdin>:1258:12
  wire [31:0] _T_131;	// <stdin>:1250:12
  wire [31:0] _T_132;	// <stdin>:1242:12
  wire [31:0] _T_133;	// <stdin>:1234:12
  wire [31:0] _T_134;	// <stdin>:1226:12
  wire [31:0] _T_135;	// <stdin>:1218:12
  wire [31:0] _T_136;	// <stdin>:1210:12
  wire [31:0] _T_137;	// <stdin>:1202:12
  wire [31:0] _T_138;	// <stdin>:1194:12
  wire [31:0] _T_139;	// <stdin>:1186:12
  wire [31:0] _T_140;	// <stdin>:1178:12
  wire [31:0] _T_141;	// <stdin>:1170:12
  wire [31:0] _T_142;	// <stdin>:1162:12
  wire [31:0] _T_143;	// <stdin>:1154:12
  wire [31:0] _T_144;	// <stdin>:1146:12
  wire [31:0] _T_145;	// <stdin>:1138:12
  wire [31:0] _T_146;	// <stdin>:1130:12
  wire [31:0] _T_147;	// <stdin>:1122:12
  wire [31:0] _T_148;	// <stdin>:1114:12
  wire [31:0] _T_149;	// <stdin>:1106:12
  wire [31:0] _T_150;	// <stdin>:1098:12
  wire [31:0] _T_151;	// <stdin>:1090:12
  wire [31:0] _T_152;	// <stdin>:1082:12
  wire [31:0] _T_153;	// <stdin>:1074:12
  wire [31:0] _T_154;	// <stdin>:1066:12
  wire [31:0] _T_155;	// <stdin>:1058:12
  wire [31:0] _T_156;	// <stdin>:1050:12
  wire [31:0] _T_157;	// <stdin>:1042:12
  wire [31:0] _T_158;	// <stdin>:1034:12
  wire [31:0] _T_159;	// <stdin>:1026:12
  wire [31:0] _T_160;	// <stdin>:1018:12
  wire [31:0] _T_161;	// <stdin>:1010:12
  wire [31:0] _T_162;	// <stdin>:1002:12
  wire [31:0] _T_163;	// <stdin>:994:12
  wire [31:0] _T_164;	// <stdin>:986:12
  wire [31:0] _T_165;	// <stdin>:978:12
  wire [31:0] _T_166;	// <stdin>:970:12
  wire [31:0] _T_167;	// <stdin>:962:12
  wire [31:0] _T_168;	// <stdin>:954:12
  wire [31:0] _T_169;	// <stdin>:946:12
  wire [31:0] _T_170;	// <stdin>:938:12
  wire [31:0] _T_171;	// <stdin>:930:12
  wire [31:0] _T_172;	// <stdin>:922:12
  wire [31:0] _T_173;	// <stdin>:914:12
  wire [31:0] _T_174;	// <stdin>:906:12
  wire [31:0] _T_175;	// <stdin>:898:12
  wire [31:0] _T_176;	// <stdin>:890:12
  wire [31:0] _T_177;	// <stdin>:882:12
  wire [31:0] _T_178;	// <stdin>:874:12
  wire [31:0] _T_179;	// <stdin>:866:12
  wire [31:0] _T_180;	// <stdin>:858:12
  wire [31:0] _T_181;	// <stdin>:850:12
  wire [31:0] _T_182;	// <stdin>:842:12
  wire [31:0] _T_183;	// <stdin>:834:12
  wire [31:0] _T_184;	// <stdin>:826:12
  wire [31:0] _T_185;	// <stdin>:818:12
  wire [31:0] _T_186;	// <stdin>:810:12
  wire [31:0] _T_187;	// <stdin>:802:12
  wire [31:0] _T_188;	// <stdin>:794:12
  wire [31:0] _T_189;	// <stdin>:786:12
  wire [31:0] _T_190;	// <stdin>:778:12
  wire [31:0] _T_191;	// <stdin>:770:12
  wire [31:0] _T_192;	// <stdin>:762:12
  wire [31:0] _T_193;	// <stdin>:754:12
  wire [31:0] _T_194;	// <stdin>:746:12
  wire [31:0] _T_195;	// <stdin>:738:12
  wire [31:0] _T_196;	// <stdin>:730:12
  wire [31:0] _T_197;	// <stdin>:722:12
  wire [31:0] _T_198;	// <stdin>:714:12
  wire [31:0] _T_199;	// <stdin>:706:12
  wire [31:0] _T_200;	// <stdin>:698:12
  wire [31:0] _T_201;	// <stdin>:690:12
  wire [31:0] _T_202;	// <stdin>:682:12
  wire [31:0] _T_203;	// <stdin>:674:12
  wire [31:0] _T_204;	// <stdin>:666:12
  wire [31:0] _T_205;	// <stdin>:658:12
  wire [31:0] _T_206;	// <stdin>:650:12
  wire [31:0] _T_207;	// <stdin>:642:12
  wire [31:0] _T_208;	// <stdin>:634:12
  wire [31:0] _T_209;	// <stdin>:626:12
  wire [31:0] _T_210;	// <stdin>:618:12
  wire [31:0] _T_211;	// <stdin>:610:12
  wire [31:0] _T_212;	// <stdin>:602:12
  wire [31:0] _T_213;	// <stdin>:594:12
  wire [31:0] _T_214;	// <stdin>:586:12
  wire [31:0] _T_215;	// <stdin>:578:12
  wire [31:0] _T_216;	// <stdin>:570:12
  wire [31:0] _T_217;	// <stdin>:562:12
  wire [31:0] _T_218;	// <stdin>:554:12
  wire [31:0] _T_219;	// <stdin>:546:12
  wire [31:0] _T_220;	// <stdin>:538:12
  wire [31:0] _T_221;	// <stdin>:530:12
  wire [31:0] _T_222;	// <stdin>:522:12
  wire [31:0] _T_223;	// <stdin>:514:12
  wire [31:0] _T_224;	// <stdin>:506:12
  wire [31:0] _T_225;	// <stdin>:498:12
  wire [31:0] _T_226;	// <stdin>:490:12
  wire [31:0] _T_227;	// <stdin>:482:12
  wire [31:0] _T_228;	// <stdin>:474:12
  wire [31:0] _T_229;	// <stdin>:466:12
  wire [31:0] _T_230;	// <stdin>:458:12
  wire [31:0] _T_231;	// <stdin>:450:12
  wire [31:0] _T_232;	// <stdin>:442:12
  wire [31:0] _T_233;	// <stdin>:434:12
  wire [31:0] _T_234;	// <stdin>:426:12
  wire [31:0] _T_235;	// <stdin>:418:12
  wire [31:0] _T_236;	// <stdin>:410:12
  wire [31:0] _T_237;	// <stdin>:402:12
  wire [31:0] _T_238;	// <stdin>:394:12
  wire [31:0] _T_239;	// <stdin>:386:12
  wire [31:0] _T_240;	// <stdin>:378:12
  wire [31:0] _T_241;	// <stdin>:370:11
  wire [31:0] _T_242;	// <stdin>:362:11
  wire [31:0] _T_243;	// <stdin>:354:11
  wire [31:0] _T_244;	// <stdin>:346:11
  wire [31:0] _T_245;	// <stdin>:338:11
  wire [31:0] _T_246;	// <stdin>:330:11
  wire [31:0] _T_247;	// <stdin>:322:11
  wire [31:0] _T_248;	// <stdin>:314:11
  wire [31:0] _T_249;	// <stdin>:306:11
  wire [31:0] _T_250;	// <stdin>:298:11
  wire [31:0] _T_251;	// <stdin>:290:11
  wire [31:0] _T_252;	// <stdin>:282:11
  wire [31:0] _T_253;	// <stdin>:274:11
  wire [31:0] _T_254;	// <stdin>:266:10
  reg  [31:0] Register_inst0;	// <stdin>:265:23
  reg  [31:0] Register_inst1;	// <stdin>:273:23
  reg  [31:0] Register_inst2;	// <stdin>:281:23
  reg  [31:0] Register_inst3;	// <stdin>:289:23
  reg  [31:0] Register_inst4;	// <stdin>:297:23
  reg  [31:0] Register_inst5;	// <stdin>:305:23
  reg  [31:0] Register_inst6;	// <stdin>:313:23
  reg  [31:0] Register_inst7;	// <stdin>:321:23
  reg  [31:0] Register_inst8;	// <stdin>:329:23
  reg  [31:0] Register_inst9;	// <stdin>:337:23
  reg  [31:0] Register_inst10;	// <stdin>:345:24
  reg  [31:0] Register_inst11;	// <stdin>:353:24
  reg  [31:0] Register_inst12;	// <stdin>:361:24
  reg  [31:0] Register_inst13;	// <stdin>:369:24
  reg  [31:0] Register_inst14;	// <stdin>:377:24
  reg  [31:0] Register_inst15;	// <stdin>:385:24
  reg  [31:0] Register_inst16;	// <stdin>:393:24
  reg  [31:0] Register_inst17;	// <stdin>:401:24
  reg  [31:0] Register_inst18;	// <stdin>:409:24
  reg  [31:0] Register_inst19;	// <stdin>:417:24
  reg  [31:0] Register_inst20;	// <stdin>:425:24
  reg  [31:0] Register_inst21;	// <stdin>:433:24
  reg  [31:0] Register_inst22;	// <stdin>:441:24
  reg  [31:0] Register_inst23;	// <stdin>:449:24
  reg  [31:0] Register_inst24;	// <stdin>:457:24
  reg  [31:0] Register_inst25;	// <stdin>:465:24
  reg  [31:0] Register_inst26;	// <stdin>:473:24
  reg  [31:0] Register_inst27;	// <stdin>:481:24
  reg  [31:0] Register_inst28;	// <stdin>:489:24
  reg  [31:0] Register_inst29;	// <stdin>:497:24
  reg  [31:0] Register_inst30;	// <stdin>:505:24
  reg  [31:0] Register_inst31;	// <stdin>:513:24
  reg  [31:0] Register_inst32;	// <stdin>:521:24
  reg  [31:0] Register_inst33;	// <stdin>:529:24
  reg  [31:0] Register_inst34;	// <stdin>:537:24
  reg  [31:0] Register_inst35;	// <stdin>:545:24
  reg  [31:0] Register_inst36;	// <stdin>:553:24
  reg  [31:0] Register_inst37;	// <stdin>:561:24
  reg  [31:0] Register_inst38;	// <stdin>:569:24
  reg  [31:0] Register_inst39;	// <stdin>:577:24
  reg  [31:0] Register_inst40;	// <stdin>:585:24
  reg  [31:0] Register_inst41;	// <stdin>:593:24
  reg  [31:0] Register_inst42;	// <stdin>:601:24
  reg  [31:0] Register_inst43;	// <stdin>:609:24
  reg  [31:0] Register_inst44;	// <stdin>:617:24
  reg  [31:0] Register_inst45;	// <stdin>:625:24
  reg  [31:0] Register_inst46;	// <stdin>:633:24
  reg  [31:0] Register_inst47;	// <stdin>:641:24
  reg  [31:0] Register_inst48;	// <stdin>:649:24
  reg  [31:0] Register_inst49;	// <stdin>:657:24
  reg  [31:0] Register_inst50;	// <stdin>:665:24
  reg  [31:0] Register_inst51;	// <stdin>:673:24
  reg  [31:0] Register_inst52;	// <stdin>:681:24
  reg  [31:0] Register_inst53;	// <stdin>:689:24
  reg  [31:0] Register_inst54;	// <stdin>:697:24
  reg  [31:0] Register_inst55;	// <stdin>:705:24
  reg  [31:0] Register_inst56;	// <stdin>:713:24
  reg  [31:0] Register_inst57;	// <stdin>:721:24
  reg  [31:0] Register_inst58;	// <stdin>:729:24
  reg  [31:0] Register_inst59;	// <stdin>:737:24
  reg  [31:0] Register_inst60;	// <stdin>:745:24
  reg  [31:0] Register_inst61;	// <stdin>:753:24
  reg  [31:0] Register_inst62;	// <stdin>:761:24
  reg  [31:0] Register_inst63;	// <stdin>:769:24
  reg  [31:0] Register_inst64;	// <stdin>:777:24
  reg  [31:0] Register_inst65;	// <stdin>:785:24
  reg  [31:0] Register_inst66;	// <stdin>:793:24
  reg  [31:0] Register_inst67;	// <stdin>:801:24
  reg  [31:0] Register_inst68;	// <stdin>:809:24
  reg  [31:0] Register_inst69;	// <stdin>:817:24
  reg  [31:0] Register_inst70;	// <stdin>:825:24
  reg  [31:0] Register_inst71;	// <stdin>:833:24
  reg  [31:0] Register_inst72;	// <stdin>:841:24
  reg  [31:0] Register_inst73;	// <stdin>:849:24
  reg  [31:0] Register_inst74;	// <stdin>:857:24
  reg  [31:0] Register_inst75;	// <stdin>:865:24
  reg  [31:0] Register_inst76;	// <stdin>:873:24
  reg  [31:0] Register_inst77;	// <stdin>:881:24
  reg  [31:0] Register_inst78;	// <stdin>:889:24
  reg  [31:0] Register_inst79;	// <stdin>:897:24
  reg  [31:0] Register_inst80;	// <stdin>:905:24
  reg  [31:0] Register_inst81;	// <stdin>:913:24
  reg  [31:0] Register_inst82;	// <stdin>:921:24
  reg  [31:0] Register_inst83;	// <stdin>:929:24
  reg  [31:0] Register_inst84;	// <stdin>:937:24
  reg  [31:0] Register_inst85;	// <stdin>:945:24
  reg  [31:0] Register_inst86;	// <stdin>:953:24
  reg  [31:0] Register_inst87;	// <stdin>:961:24
  reg  [31:0] Register_inst88;	// <stdin>:969:24
  reg  [31:0] Register_inst89;	// <stdin>:977:24
  reg  [31:0] Register_inst90;	// <stdin>:985:24
  reg  [31:0] Register_inst91;	// <stdin>:993:24
  reg  [31:0] Register_inst92;	// <stdin>:1001:24
  reg  [31:0] Register_inst93;	// <stdin>:1009:24
  reg  [31:0] Register_inst94;	// <stdin>:1017:24
  reg  [31:0] Register_inst95;	// <stdin>:1025:24
  reg  [31:0] Register_inst96;	// <stdin>:1033:24
  reg  [31:0] Register_inst97;	// <stdin>:1041:24
  reg  [31:0] Register_inst98;	// <stdin>:1049:24
  reg  [31:0] Register_inst99;	// <stdin>:1057:24
  reg  [31:0] Register_inst100;	// <stdin>:1065:25
  reg  [31:0] Register_inst101;	// <stdin>:1073:25
  reg  [31:0] Register_inst102;	// <stdin>:1081:25
  reg  [31:0] Register_inst103;	// <stdin>:1089:25
  reg  [31:0] Register_inst104;	// <stdin>:1097:25
  reg  [31:0] Register_inst105;	// <stdin>:1105:25
  reg  [31:0] Register_inst106;	// <stdin>:1113:25
  reg  [31:0] Register_inst107;	// <stdin>:1121:25
  reg  [31:0] Register_inst108;	// <stdin>:1129:25
  reg  [31:0] Register_inst109;	// <stdin>:1137:25
  reg  [31:0] Register_inst110;	// <stdin>:1145:25
  reg  [31:0] Register_inst111;	// <stdin>:1153:25
  reg  [31:0] Register_inst112;	// <stdin>:1161:25
  reg  [31:0] Register_inst113;	// <stdin>:1169:25
  reg  [31:0] Register_inst114;	// <stdin>:1177:25
  reg  [31:0] Register_inst115;	// <stdin>:1185:25
  reg  [31:0] Register_inst116;	// <stdin>:1193:25
  reg  [31:0] Register_inst117;	// <stdin>:1201:25
  reg  [31:0] Register_inst118;	// <stdin>:1209:25
  reg  [31:0] Register_inst119;	// <stdin>:1217:25
  reg  [31:0] Register_inst120;	// <stdin>:1225:25
  reg  [31:0] Register_inst121;	// <stdin>:1233:25
  reg  [31:0] Register_inst122;	// <stdin>:1241:25
  reg  [31:0] Register_inst123;	// <stdin>:1249:25
  reg  [31:0] Register_inst124;	// <stdin>:1257:25
  reg  [31:0] Register_inst125;	// <stdin>:1265:25
  reg  [31:0] Register_inst126;	// <stdin>:1273:25
  reg  [31:0] Register_inst127;	// <stdin>:1281:25
  reg  [31:0] Register_inst128;	// <stdin>:1289:25
  reg  [31:0] Register_inst129;	// <stdin>:1297:25
  reg  [31:0] Register_inst130;	// <stdin>:1305:25
  reg  [31:0] Register_inst131;	// <stdin>:1313:25
  reg  [31:0] Register_inst132;	// <stdin>:1321:25
  reg  [31:0] Register_inst133;	// <stdin>:1329:25
  reg  [31:0] Register_inst134;	// <stdin>:1337:25
  reg  [31:0] Register_inst135;	// <stdin>:1345:25
  reg  [31:0] Register_inst136;	// <stdin>:1353:25
  reg  [31:0] Register_inst137;	// <stdin>:1361:25
  reg  [31:0] Register_inst138;	// <stdin>:1369:25
  reg  [31:0] Register_inst139;	// <stdin>:1377:25
  reg  [31:0] Register_inst140;	// <stdin>:1385:25
  reg  [31:0] Register_inst141;	// <stdin>:1393:25
  reg  [31:0] Register_inst142;	// <stdin>:1401:25
  reg  [31:0] Register_inst143;	// <stdin>:1409:25
  reg  [31:0] Register_inst144;	// <stdin>:1417:25
  reg  [31:0] Register_inst145;	// <stdin>:1425:25
  reg  [31:0] Register_inst146;	// <stdin>:1433:25
  reg  [31:0] Register_inst147;	// <stdin>:1441:25
  reg  [31:0] Register_inst148;	// <stdin>:1449:25
  reg  [31:0] Register_inst149;	// <stdin>:1457:25
  reg  [31:0] Register_inst150;	// <stdin>:1465:25
  reg  [31:0] Register_inst151;	// <stdin>:1473:25
  reg  [31:0] Register_inst152;	// <stdin>:1481:25
  reg  [31:0] Register_inst153;	// <stdin>:1489:25
  reg  [31:0] Register_inst154;	// <stdin>:1497:25
  reg  [31:0] Register_inst155;	// <stdin>:1505:25
  reg  [31:0] Register_inst156;	// <stdin>:1513:25
  reg  [31:0] Register_inst157;	// <stdin>:1521:25
  reg  [31:0] Register_inst158;	// <stdin>:1529:25
  reg  [31:0] Register_inst159;	// <stdin>:1537:25
  reg  [31:0] Register_inst160;	// <stdin>:1545:25
  reg  [31:0] Register_inst161;	// <stdin>:1553:25
  reg  [31:0] Register_inst162;	// <stdin>:1561:25
  reg  [31:0] Register_inst163;	// <stdin>:1569:25
  reg  [31:0] Register_inst164;	// <stdin>:1577:25
  reg  [31:0] Register_inst165;	// <stdin>:1585:25
  reg  [31:0] Register_inst166;	// <stdin>:1593:25
  reg  [31:0] Register_inst167;	// <stdin>:1601:25
  reg  [31:0] Register_inst168;	// <stdin>:1609:25
  reg  [31:0] Register_inst169;	// <stdin>:1617:25
  reg  [31:0] Register_inst170;	// <stdin>:1625:25
  reg  [31:0] Register_inst171;	// <stdin>:1633:25
  reg  [31:0] Register_inst172;	// <stdin>:1641:25
  reg  [31:0] Register_inst173;	// <stdin>:1649:25
  reg  [31:0] Register_inst174;	// <stdin>:1657:25
  reg  [31:0] Register_inst175;	// <stdin>:1665:25
  reg  [31:0] Register_inst176;	// <stdin>:1673:25
  reg  [31:0] Register_inst177;	// <stdin>:1681:25
  reg  [31:0] Register_inst178;	// <stdin>:1689:25
  reg  [31:0] Register_inst179;	// <stdin>:1697:25
  reg  [31:0] Register_inst180;	// <stdin>:1705:25
  reg  [31:0] Register_inst181;	// <stdin>:1713:25
  reg  [31:0] Register_inst182;	// <stdin>:1721:25
  reg  [31:0] Register_inst183;	// <stdin>:1729:25
  reg  [31:0] Register_inst184;	// <stdin>:1737:25
  reg  [31:0] Register_inst185;	// <stdin>:1745:25
  reg  [31:0] Register_inst186;	// <stdin>:1753:25
  reg  [31:0] Register_inst187;	// <stdin>:1761:25
  reg  [31:0] Register_inst188;	// <stdin>:1769:25
  reg  [31:0] Register_inst189;	// <stdin>:1777:25
  reg  [31:0] Register_inst190;	// <stdin>:1785:25
  reg  [31:0] Register_inst191;	// <stdin>:1793:25
  reg  [31:0] Register_inst192;	// <stdin>:1801:25
  reg  [31:0] Register_inst193;	// <stdin>:1809:25
  reg  [31:0] Register_inst194;	// <stdin>:1817:25
  reg  [31:0] Register_inst195;	// <stdin>:1825:25
  reg  [31:0] Register_inst196;	// <stdin>:1833:25
  reg  [31:0] Register_inst197;	// <stdin>:1841:25
  reg  [31:0] Register_inst198;	// <stdin>:1849:25
  reg  [31:0] Register_inst199;	// <stdin>:1857:25
  reg  [31:0] Register_inst200;	// <stdin>:1865:25
  reg  [31:0] Register_inst201;	// <stdin>:1873:25
  reg  [31:0] Register_inst202;	// <stdin>:1881:25
  reg  [31:0] Register_inst203;	// <stdin>:1889:25
  reg  [31:0] Register_inst204;	// <stdin>:1897:25
  reg  [31:0] Register_inst205;	// <stdin>:1905:25
  reg  [31:0] Register_inst206;	// <stdin>:1913:25
  reg  [31:0] Register_inst207;	// <stdin>:1921:25
  reg  [31:0] Register_inst208;	// <stdin>:1929:25
  reg  [31:0] Register_inst209;	// <stdin>:1937:25
  reg  [31:0] Register_inst210;	// <stdin>:1945:25
  reg  [31:0] Register_inst211;	// <stdin>:1953:25
  reg  [31:0] Register_inst212;	// <stdin>:1961:25
  reg  [31:0] Register_inst213;	// <stdin>:1969:25
  reg  [31:0] Register_inst214;	// <stdin>:1977:25
  reg  [31:0] Register_inst215;	// <stdin>:1985:25
  reg  [31:0] Register_inst216;	// <stdin>:1993:25
  reg  [31:0] Register_inst217;	// <stdin>:2001:25
  reg  [31:0] Register_inst218;	// <stdin>:2009:25
  reg  [31:0] Register_inst219;	// <stdin>:2017:25
  reg  [31:0] Register_inst220;	// <stdin>:2025:25
  reg  [31:0] Register_inst221;	// <stdin>:2033:25
  reg  [31:0] Register_inst222;	// <stdin>:2041:25
  reg  [31:0] Register_inst223;	// <stdin>:2049:25
  reg  [31:0] Register_inst224;	// <stdin>:2057:25
  reg  [31:0] Register_inst225;	// <stdin>:2065:25
  reg  [31:0] Register_inst226;	// <stdin>:2073:25
  reg  [31:0] Register_inst227;	// <stdin>:2081:25
  reg  [31:0] Register_inst228;	// <stdin>:2089:25
  reg  [31:0] Register_inst229;	// <stdin>:2097:25
  reg  [31:0] Register_inst230;	// <stdin>:2105:25
  reg  [31:0] Register_inst231;	// <stdin>:2113:25
  reg  [31:0] Register_inst232;	// <stdin>:2121:25
  reg  [31:0] Register_inst233;	// <stdin>:2129:25
  reg  [31:0] Register_inst234;	// <stdin>:2137:25
  reg  [31:0] Register_inst235;	// <stdin>:2145:25
  reg  [31:0] Register_inst236;	// <stdin>:2153:25
  reg  [31:0] Register_inst237;	// <stdin>:2161:25
  reg  [31:0] Register_inst238;	// <stdin>:2169:25
  reg  [31:0] Register_inst239;	// <stdin>:2177:25
  reg  [31:0] Register_inst240;	// <stdin>:2185:25
  reg  [31:0] Register_inst241;	// <stdin>:2193:25
  reg  [31:0] Register_inst242;	// <stdin>:2201:25
  reg  [31:0] Register_inst243;	// <stdin>:2209:25
  reg  [31:0] Register_inst244;	// <stdin>:2217:25
  reg  [31:0] Register_inst245;	// <stdin>:2225:25
  reg  [31:0] Register_inst246;	// <stdin>:2233:25
  reg  [31:0] Register_inst247;	// <stdin>:2241:25
  reg  [31:0] Register_inst248;	// <stdin>:2249:25
  reg  [31:0] Register_inst249;	// <stdin>:2257:25
  reg  [31:0] Register_inst250;	// <stdin>:2265:25
  reg  [31:0] Register_inst251;	// <stdin>:2273:25
  reg  [31:0] Register_inst252;	// <stdin>:2281:25
  reg  [31:0] Register_inst253;	// <stdin>:2289:25
  reg  [31:0] Register_inst254;	// <stdin>:2297:25
  reg  [31:0] Register_inst255;	// <stdin>:2305:25

  wire [31:0] _T_255 = ({{_T_254}, {write_0.data}})[write_0.addr == 8'h0 & write_0_en];	// <stdin>:258:14, :259:10, :260:10, :261:10, :262:10, :263:10, :264:10, :266:10
  assign _T_254 = Register_inst0;	// <stdin>:266:10
  wire [31:0] _T_256 = ({{_T_253}, {write_0.data}})[write_0.addr == 8'h1 & write_0_en];	// <stdin>:257:14, :267:10, :268:10, :269:10, :270:11, :271:11, :272:11, :274:11
  assign _T_253 = Register_inst1;	// <stdin>:274:11
  wire [31:0] _T_257 = ({{_T_252}, {write_0.data}})[write_0.addr == 8'h2 & write_0_en];	// <stdin>:256:14, :275:11, :276:11, :277:11, :278:11, :279:11, :280:11, :282:11
  assign _T_252 = Register_inst2;	// <stdin>:282:11
  wire [31:0] _T_258 = ({{_T_251}, {write_0.data}})[write_0.addr == 8'h3 & write_0_en];	// <stdin>:255:14, :283:11, :284:11, :285:11, :286:11, :287:11, :288:11, :290:11
  assign _T_251 = Register_inst3;	// <stdin>:290:11
  wire [31:0] _T_259 = ({{_T_250}, {write_0.data}})[write_0.addr == 8'h4 & write_0_en];	// <stdin>:254:14, :291:11, :292:11, :293:11, :294:11, :295:11, :296:11, :298:11
  assign _T_250 = Register_inst4;	// <stdin>:298:11
  wire [31:0] _T_260 = ({{_T_249}, {write_0.data}})[write_0.addr == 8'h5 & write_0_en];	// <stdin>:253:14, :299:11, :300:11, :301:11, :302:11, :303:11, :304:11, :306:11
  assign _T_249 = Register_inst5;	// <stdin>:306:11
  wire [31:0] _T_261 = ({{_T_248}, {write_0.data}})[write_0.addr == 8'h6 & write_0_en];	// <stdin>:252:14, :307:11, :308:11, :309:11, :310:11, :311:11, :312:11, :314:11
  assign _T_248 = Register_inst6;	// <stdin>:314:11
  wire [31:0] _T_262 = ({{_T_247}, {write_0.data}})[write_0.addr == 8'h7 & write_0_en];	// <stdin>:251:14, :315:11, :316:11, :317:11, :318:11, :319:11, :320:11, :322:11
  assign _T_247 = Register_inst7;	// <stdin>:322:11
  wire [31:0] _T_263 = ({{_T_246}, {write_0.data}})[write_0.addr == 8'h8 & write_0_en];	// <stdin>:250:14, :323:11, :324:11, :325:11, :326:11, :327:11, :328:11, :330:11
  assign _T_246 = Register_inst8;	// <stdin>:330:11
  wire [31:0] _T_264 = ({{_T_245}, {write_0.data}})[write_0.addr == 8'h9 & write_0_en];	// <stdin>:249:14, :331:11, :332:11, :333:11, :334:11, :335:11, :336:11, :338:11
  assign _T_245 = Register_inst9;	// <stdin>:338:11
  wire [31:0] _T_265 = ({{_T_244}, {write_0.data}})[write_0.addr == 8'hA & write_0_en];	// <stdin>:248:15, :339:11, :340:11, :341:11, :342:11, :343:11, :344:11, :346:11
  assign _T_244 = Register_inst10;	// <stdin>:346:11
  wire [31:0] _T_266 = ({{_T_243}, {write_0.data}})[write_0.addr == 8'hB & write_0_en];	// <stdin>:247:15, :347:11, :348:11, :349:11, :350:11, :351:11, :352:11, :354:11
  assign _T_243 = Register_inst11;	// <stdin>:354:11
  wire [31:0] _T_267 = ({{_T_242}, {write_0.data}})[write_0.addr == 8'hC & write_0_en];	// <stdin>:246:15, :355:11, :356:11, :357:11, :358:11, :359:11, :360:11, :362:11
  assign _T_242 = Register_inst12;	// <stdin>:362:11
  wire [31:0] _T_268 = ({{_T_241}, {write_0.data}})[write_0.addr == 8'hD & write_0_en];	// <stdin>:245:15, :363:11, :364:11, :365:11, :366:11, :367:11, :368:11, :370:11
  assign _T_241 = Register_inst13;	// <stdin>:370:11
  wire [31:0] _T_269 = ({{_T_240}, {write_0.data}})[write_0.addr == 8'hE & write_0_en];	// <stdin>:244:15, :371:11, :372:11, :373:12, :374:12, :375:12, :376:12, :378:12
  assign _T_240 = Register_inst14;	// <stdin>:378:12
  wire [31:0] _T_270 = ({{_T_239}, {write_0.data}})[write_0.addr == 8'hF & write_0_en];	// <stdin>:243:15, :379:12, :380:12, :381:12, :382:12, :383:12, :384:12, :386:12
  assign _T_239 = Register_inst15;	// <stdin>:386:12
  wire [31:0] _T_271 = ({{_T_238}, {write_0.data}})[write_0.addr == 8'h10 & write_0_en];	// <stdin>:242:15, :387:12, :388:12, :389:12, :390:12, :391:12, :392:12, :394:12
  assign _T_238 = Register_inst16;	// <stdin>:394:12
  wire [31:0] _T_272 = ({{_T_237}, {write_0.data}})[write_0.addr == 8'h11 & write_0_en];	// <stdin>:241:15, :395:12, :396:12, :397:12, :398:12, :399:12, :400:12, :402:12
  assign _T_237 = Register_inst17;	// <stdin>:402:12
  wire [31:0] _T_273 = ({{_T_236}, {write_0.data}})[write_0.addr == 8'h12 & write_0_en];	// <stdin>:240:15, :403:12, :404:12, :405:12, :406:12, :407:12, :408:12, :410:12
  assign _T_236 = Register_inst18;	// <stdin>:410:12
  wire [31:0] _T_274 = ({{_T_235}, {write_0.data}})[write_0.addr == 8'h13 & write_0_en];	// <stdin>:239:15, :411:12, :412:12, :413:12, :414:12, :415:12, :416:12, :418:12
  assign _T_235 = Register_inst19;	// <stdin>:418:12
  wire [31:0] _T_275 = ({{_T_234}, {write_0.data}})[write_0.addr == 8'h14 & write_0_en];	// <stdin>:238:15, :419:12, :420:12, :421:12, :422:12, :423:12, :424:12, :426:12
  assign _T_234 = Register_inst20;	// <stdin>:426:12
  wire [31:0] _T_276 = ({{_T_233}, {write_0.data}})[write_0.addr == 8'h15 & write_0_en];	// <stdin>:237:15, :427:12, :428:12, :429:12, :430:12, :431:12, :432:12, :434:12
  assign _T_233 = Register_inst21;	// <stdin>:434:12
  wire [31:0] _T_277 = ({{_T_232}, {write_0.data}})[write_0.addr == 8'h16 & write_0_en];	// <stdin>:236:15, :435:12, :436:12, :437:12, :438:12, :439:12, :440:12, :442:12
  assign _T_232 = Register_inst22;	// <stdin>:442:12
  wire [31:0] _T_278 = ({{_T_231}, {write_0.data}})[write_0.addr == 8'h17 & write_0_en];	// <stdin>:235:15, :443:12, :444:12, :445:12, :446:12, :447:12, :448:12, :450:12
  assign _T_231 = Register_inst23;	// <stdin>:450:12
  wire [31:0] _T_279 = ({{_T_230}, {write_0.data}})[write_0.addr == 8'h18 & write_0_en];	// <stdin>:234:15, :451:12, :452:12, :453:12, :454:12, :455:12, :456:12, :458:12
  assign _T_230 = Register_inst24;	// <stdin>:458:12
  wire [31:0] _T_280 = ({{_T_229}, {write_0.data}})[write_0.addr == 8'h19 & write_0_en];	// <stdin>:233:15, :459:12, :460:12, :461:12, :462:12, :463:12, :464:12, :466:12
  assign _T_229 = Register_inst25;	// <stdin>:466:12
  wire [31:0] _T_281 = ({{_T_228}, {write_0.data}})[write_0.addr == 8'h1A & write_0_en];	// <stdin>:232:15, :467:12, :468:12, :469:12, :470:12, :471:12, :472:12, :474:12
  assign _T_228 = Register_inst26;	// <stdin>:474:12
  wire [31:0] _T_282 = ({{_T_227}, {write_0.data}})[write_0.addr == 8'h1B & write_0_en];	// <stdin>:231:15, :475:12, :476:12, :477:12, :478:12, :479:12, :480:12, :482:12
  assign _T_227 = Register_inst27;	// <stdin>:482:12
  wire [31:0] _T_283 = ({{_T_226}, {write_0.data}})[write_0.addr == 8'h1C & write_0_en];	// <stdin>:230:15, :483:12, :484:12, :485:12, :486:12, :487:12, :488:12, :490:12
  assign _T_226 = Register_inst28;	// <stdin>:490:12
  wire [31:0] _T_284 = ({{_T_225}, {write_0.data}})[write_0.addr == 8'h1D & write_0_en];	// <stdin>:229:15, :491:12, :492:12, :493:12, :494:12, :495:12, :496:12, :498:12
  assign _T_225 = Register_inst29;	// <stdin>:498:12
  wire [31:0] _T_285 = ({{_T_224}, {write_0.data}})[write_0.addr == 8'h1E & write_0_en];	// <stdin>:228:15, :499:12, :500:12, :501:12, :502:12, :503:12, :504:12, :506:12
  assign _T_224 = Register_inst30;	// <stdin>:506:12
  wire [31:0] _T_286 = ({{_T_223}, {write_0.data}})[write_0.addr == 8'h1F & write_0_en];	// <stdin>:227:15, :507:12, :508:12, :509:12, :510:12, :511:12, :512:12, :514:12
  assign _T_223 = Register_inst31;	// <stdin>:514:12
  wire [31:0] _T_287 = ({{_T_222}, {write_0.data}})[write_0.addr == 8'h20 & write_0_en];	// <stdin>:226:15, :515:12, :516:12, :517:12, :518:12, :519:12, :520:12, :522:12
  assign _T_222 = Register_inst32;	// <stdin>:522:12
  wire [31:0] _T_288 = ({{_T_221}, {write_0.data}})[write_0.addr == 8'h21 & write_0_en];	// <stdin>:225:15, :523:12, :524:12, :525:12, :526:12, :527:12, :528:12, :530:12
  assign _T_221 = Register_inst33;	// <stdin>:530:12
  wire [31:0] _T_289 = ({{_T_220}, {write_0.data}})[write_0.addr == 8'h22 & write_0_en];	// <stdin>:224:15, :531:12, :532:12, :533:12, :534:12, :535:12, :536:12, :538:12
  assign _T_220 = Register_inst34;	// <stdin>:538:12
  wire [31:0] _T_290 = ({{_T_219}, {write_0.data}})[write_0.addr == 8'h23 & write_0_en];	// <stdin>:223:15, :539:12, :540:12, :541:12, :542:12, :543:12, :544:12, :546:12
  assign _T_219 = Register_inst35;	// <stdin>:546:12
  wire [31:0] _T_291 = ({{_T_218}, {write_0.data}})[write_0.addr == 8'h24 & write_0_en];	// <stdin>:222:15, :547:12, :548:12, :549:12, :550:12, :551:12, :552:12, :554:12
  assign _T_218 = Register_inst36;	// <stdin>:554:12
  wire [31:0] _T_292 = ({{_T_217}, {write_0.data}})[write_0.addr == 8'h25 & write_0_en];	// <stdin>:221:15, :555:12, :556:12, :557:12, :558:12, :559:12, :560:12, :562:12
  assign _T_217 = Register_inst37;	// <stdin>:562:12
  wire [31:0] _T_293 = ({{_T_216}, {write_0.data}})[write_0.addr == 8'h26 & write_0_en];	// <stdin>:220:15, :563:12, :564:12, :565:12, :566:12, :567:12, :568:12, :570:12
  assign _T_216 = Register_inst38;	// <stdin>:570:12
  wire [31:0] _T_294 = ({{_T_215}, {write_0.data}})[write_0.addr == 8'h27 & write_0_en];	// <stdin>:219:15, :571:12, :572:12, :573:12, :574:12, :575:12, :576:12, :578:12
  assign _T_215 = Register_inst39;	// <stdin>:578:12
  wire [31:0] _T_295 = ({{_T_214}, {write_0.data}})[write_0.addr == 8'h28 & write_0_en];	// <stdin>:218:15, :579:12, :580:12, :581:12, :582:12, :583:12, :584:12, :586:12
  assign _T_214 = Register_inst40;	// <stdin>:586:12
  wire [31:0] _T_296 = ({{_T_213}, {write_0.data}})[write_0.addr == 8'h29 & write_0_en];	// <stdin>:217:15, :587:12, :588:12, :589:12, :590:12, :591:12, :592:12, :594:12
  assign _T_213 = Register_inst41;	// <stdin>:594:12
  wire [31:0] _T_297 = ({{_T_212}, {write_0.data}})[write_0.addr == 8'h2A & write_0_en];	// <stdin>:216:15, :595:12, :596:12, :597:12, :598:12, :599:12, :600:12, :602:12
  assign _T_212 = Register_inst42;	// <stdin>:602:12
  wire [31:0] _T_298 = ({{_T_211}, {write_0.data}})[write_0.addr == 8'h2B & write_0_en];	// <stdin>:215:15, :603:12, :604:12, :605:12, :606:12, :607:12, :608:12, :610:12
  assign _T_211 = Register_inst43;	// <stdin>:610:12
  wire [31:0] _T_299 = ({{_T_210}, {write_0.data}})[write_0.addr == 8'h2C & write_0_en];	// <stdin>:214:15, :611:12, :612:12, :613:12, :614:12, :615:12, :616:12, :618:12
  assign _T_210 = Register_inst44;	// <stdin>:618:12
  wire [31:0] _T_300 = ({{_T_209}, {write_0.data}})[write_0.addr == 8'h2D & write_0_en];	// <stdin>:213:15, :619:12, :620:12, :621:12, :622:12, :623:12, :624:12, :626:12
  assign _T_209 = Register_inst45;	// <stdin>:626:12
  wire [31:0] _T_301 = ({{_T_208}, {write_0.data}})[write_0.addr == 8'h2E & write_0_en];	// <stdin>:212:15, :627:12, :628:12, :629:12, :630:12, :631:12, :632:12, :634:12
  assign _T_208 = Register_inst46;	// <stdin>:634:12
  wire [31:0] _T_302 = ({{_T_207}, {write_0.data}})[write_0.addr == 8'h2F & write_0_en];	// <stdin>:211:15, :635:12, :636:12, :637:12, :638:12, :639:12, :640:12, :642:12
  assign _T_207 = Register_inst47;	// <stdin>:642:12
  wire [31:0] _T_303 = ({{_T_206}, {write_0.data}})[write_0.addr == 8'h30 & write_0_en];	// <stdin>:210:15, :643:12, :644:12, :645:12, :646:12, :647:12, :648:12, :650:12
  assign _T_206 = Register_inst48;	// <stdin>:650:12
  wire [31:0] _T_304 = ({{_T_205}, {write_0.data}})[write_0.addr == 8'h31 & write_0_en];	// <stdin>:209:15, :651:12, :652:12, :653:12, :654:12, :655:12, :656:12, :658:12
  assign _T_205 = Register_inst49;	// <stdin>:658:12
  wire [31:0] _T_305 = ({{_T_204}, {write_0.data}})[write_0.addr == 8'h32 & write_0_en];	// <stdin>:208:15, :659:12, :660:12, :661:12, :662:12, :663:12, :664:12, :666:12
  assign _T_204 = Register_inst50;	// <stdin>:666:12
  wire [31:0] _T_306 = ({{_T_203}, {write_0.data}})[write_0.addr == 8'h33 & write_0_en];	// <stdin>:207:15, :667:12, :668:12, :669:12, :670:12, :671:12, :672:12, :674:12
  assign _T_203 = Register_inst51;	// <stdin>:674:12
  wire [31:0] _T_307 = ({{_T_202}, {write_0.data}})[write_0.addr == 8'h34 & write_0_en];	// <stdin>:206:15, :675:12, :676:12, :677:12, :678:12, :679:12, :680:12, :682:12
  assign _T_202 = Register_inst52;	// <stdin>:682:12
  wire [31:0] _T_308 = ({{_T_201}, {write_0.data}})[write_0.addr == 8'h35 & write_0_en];	// <stdin>:205:15, :683:12, :684:12, :685:12, :686:12, :687:12, :688:12, :690:12
  assign _T_201 = Register_inst53;	// <stdin>:690:12
  wire [31:0] _T_309 = ({{_T_200}, {write_0.data}})[write_0.addr == 8'h36 & write_0_en];	// <stdin>:204:15, :691:12, :692:12, :693:12, :694:12, :695:12, :696:12, :698:12
  assign _T_200 = Register_inst54;	// <stdin>:698:12
  wire [31:0] _T_310 = ({{_T_199}, {write_0.data}})[write_0.addr == 8'h37 & write_0_en];	// <stdin>:203:15, :699:12, :700:12, :701:12, :702:12, :703:12, :704:12, :706:12
  assign _T_199 = Register_inst55;	// <stdin>:706:12
  wire [31:0] _T_311 = ({{_T_198}, {write_0.data}})[write_0.addr == 8'h38 & write_0_en];	// <stdin>:202:15, :707:12, :708:12, :709:12, :710:12, :711:12, :712:12, :714:12
  assign _T_198 = Register_inst56;	// <stdin>:714:12
  wire [31:0] _T_312 = ({{_T_197}, {write_0.data}})[write_0.addr == 8'h39 & write_0_en];	// <stdin>:201:15, :715:12, :716:12, :717:12, :718:12, :719:12, :720:12, :722:12
  assign _T_197 = Register_inst57;	// <stdin>:722:12
  wire [31:0] _T_313 = ({{_T_196}, {write_0.data}})[write_0.addr == 8'h3A & write_0_en];	// <stdin>:200:15, :723:12, :724:12, :725:12, :726:12, :727:12, :728:12, :730:12
  assign _T_196 = Register_inst58;	// <stdin>:730:12
  wire [31:0] _T_314 = ({{_T_195}, {write_0.data}})[write_0.addr == 8'h3B & write_0_en];	// <stdin>:199:15, :731:12, :732:12, :733:12, :734:12, :735:12, :736:12, :738:12
  assign _T_195 = Register_inst59;	// <stdin>:738:12
  wire [31:0] _T_315 = ({{_T_194}, {write_0.data}})[write_0.addr == 8'h3C & write_0_en];	// <stdin>:198:15, :739:12, :740:12, :741:12, :742:12, :743:12, :744:12, :746:12
  assign _T_194 = Register_inst60;	// <stdin>:746:12
  wire [31:0] _T_316 = ({{_T_193}, {write_0.data}})[write_0.addr == 8'h3D & write_0_en];	// <stdin>:197:15, :747:12, :748:12, :749:12, :750:12, :751:12, :752:12, :754:12
  assign _T_193 = Register_inst61;	// <stdin>:754:12
  wire [31:0] _T_317 = ({{_T_192}, {write_0.data}})[write_0.addr == 8'h3E & write_0_en];	// <stdin>:196:15, :755:12, :756:12, :757:12, :758:12, :759:12, :760:12, :762:12
  assign _T_192 = Register_inst62;	// <stdin>:762:12
  wire [31:0] _T_318 = ({{_T_191}, {write_0.data}})[write_0.addr == 8'h3F & write_0_en];	// <stdin>:195:15, :763:12, :764:12, :765:12, :766:12, :767:12, :768:12, :770:12
  assign _T_191 = Register_inst63;	// <stdin>:770:12
  wire [31:0] _T_319 = ({{_T_190}, {write_0.data}})[write_0.addr == 8'h40 & write_0_en];	// <stdin>:194:15, :771:12, :772:12, :773:12, :774:12, :775:12, :776:12, :778:12
  assign _T_190 = Register_inst64;	// <stdin>:778:12
  wire [31:0] _T_320 = ({{_T_189}, {write_0.data}})[write_0.addr == 8'h41 & write_0_en];	// <stdin>:193:15, :779:12, :780:12, :781:12, :782:12, :783:12, :784:12, :786:12
  assign _T_189 = Register_inst65;	// <stdin>:786:12
  wire [31:0] _T_321 = ({{_T_188}, {write_0.data}})[write_0.addr == 8'h42 & write_0_en];	// <stdin>:192:15, :787:12, :788:12, :789:12, :790:12, :791:12, :792:12, :794:12
  assign _T_188 = Register_inst66;	// <stdin>:794:12
  wire [31:0] _T_322 = ({{_T_187}, {write_0.data}})[write_0.addr == 8'h43 & write_0_en];	// <stdin>:191:15, :795:12, :796:12, :797:12, :798:12, :799:12, :800:12, :802:12
  assign _T_187 = Register_inst67;	// <stdin>:802:12
  wire [31:0] _T_323 = ({{_T_186}, {write_0.data}})[write_0.addr == 8'h44 & write_0_en];	// <stdin>:190:15, :803:12, :804:12, :805:12, :806:12, :807:12, :808:12, :810:12
  assign _T_186 = Register_inst68;	// <stdin>:810:12
  wire [31:0] _T_324 = ({{_T_185}, {write_0.data}})[write_0.addr == 8'h45 & write_0_en];	// <stdin>:189:15, :811:12, :812:12, :813:12, :814:12, :815:12, :816:12, :818:12
  assign _T_185 = Register_inst69;	// <stdin>:818:12
  wire [31:0] _T_325 = ({{_T_184}, {write_0.data}})[write_0.addr == 8'h46 & write_0_en];	// <stdin>:188:15, :819:12, :820:12, :821:12, :822:12, :823:12, :824:12, :826:12
  assign _T_184 = Register_inst70;	// <stdin>:826:12
  wire [31:0] _T_326 = ({{_T_183}, {write_0.data}})[write_0.addr == 8'h47 & write_0_en];	// <stdin>:187:15, :827:12, :828:12, :829:12, :830:12, :831:12, :832:12, :834:12
  assign _T_183 = Register_inst71;	// <stdin>:834:12
  wire [31:0] _T_327 = ({{_T_182}, {write_0.data}})[write_0.addr == 8'h48 & write_0_en];	// <stdin>:186:15, :835:12, :836:12, :837:12, :838:12, :839:12, :840:12, :842:12
  assign _T_182 = Register_inst72;	// <stdin>:842:12
  wire [31:0] _T_328 = ({{_T_181}, {write_0.data}})[write_0.addr == 8'h49 & write_0_en];	// <stdin>:185:15, :843:12, :844:12, :845:12, :846:12, :847:12, :848:12, :850:12
  assign _T_181 = Register_inst73;	// <stdin>:850:12
  wire [31:0] _T_329 = ({{_T_180}, {write_0.data}})[write_0.addr == 8'h4A & write_0_en];	// <stdin>:184:15, :851:12, :852:12, :853:12, :854:12, :855:12, :856:12, :858:12
  assign _T_180 = Register_inst74;	// <stdin>:858:12
  wire [31:0] _T_330 = ({{_T_179}, {write_0.data}})[write_0.addr == 8'h4B & write_0_en];	// <stdin>:183:15, :859:12, :860:12, :861:12, :862:12, :863:12, :864:12, :866:12
  assign _T_179 = Register_inst75;	// <stdin>:866:12
  wire [31:0] _T_331 = ({{_T_178}, {write_0.data}})[write_0.addr == 8'h4C & write_0_en];	// <stdin>:182:15, :867:12, :868:12, :869:12, :870:12, :871:12, :872:12, :874:12
  assign _T_178 = Register_inst76;	// <stdin>:874:12
  wire [31:0] _T_332 = ({{_T_177}, {write_0.data}})[write_0.addr == 8'h4D & write_0_en];	// <stdin>:181:15, :875:12, :876:12, :877:12, :878:12, :879:12, :880:12, :882:12
  assign _T_177 = Register_inst77;	// <stdin>:882:12
  wire [31:0] _T_333 = ({{_T_176}, {write_0.data}})[write_0.addr == 8'h4E & write_0_en];	// <stdin>:180:15, :883:12, :884:12, :885:12, :886:12, :887:12, :888:12, :890:12
  assign _T_176 = Register_inst78;	// <stdin>:890:12
  wire [31:0] _T_334 = ({{_T_175}, {write_0.data}})[write_0.addr == 8'h4F & write_0_en];	// <stdin>:179:15, :891:12, :892:12, :893:12, :894:12, :895:12, :896:12, :898:12
  assign _T_175 = Register_inst79;	// <stdin>:898:12
  wire [31:0] _T_335 = ({{_T_174}, {write_0.data}})[write_0.addr == 8'h50 & write_0_en];	// <stdin>:178:15, :899:12, :900:12, :901:12, :902:12, :903:12, :904:12, :906:12
  assign _T_174 = Register_inst80;	// <stdin>:906:12
  wire [31:0] _T_336 = ({{_T_173}, {write_0.data}})[write_0.addr == 8'h51 & write_0_en];	// <stdin>:177:15, :907:12, :908:12, :909:12, :910:12, :911:12, :912:12, :914:12
  assign _T_173 = Register_inst81;	// <stdin>:914:12
  wire [31:0] _T_337 = ({{_T_172}, {write_0.data}})[write_0.addr == 8'h52 & write_0_en];	// <stdin>:176:15, :915:12, :916:12, :917:12, :918:12, :919:12, :920:12, :922:12
  assign _T_172 = Register_inst82;	// <stdin>:922:12
  wire [31:0] _T_338 = ({{_T_171}, {write_0.data}})[write_0.addr == 8'h53 & write_0_en];	// <stdin>:175:15, :923:12, :924:12, :925:12, :926:12, :927:12, :928:12, :930:12
  assign _T_171 = Register_inst83;	// <stdin>:930:12
  wire [31:0] _T_339 = ({{_T_170}, {write_0.data}})[write_0.addr == 8'h54 & write_0_en];	// <stdin>:174:15, :931:12, :932:12, :933:12, :934:12, :935:12, :936:12, :938:12
  assign _T_170 = Register_inst84;	// <stdin>:938:12
  wire [31:0] _T_340 = ({{_T_169}, {write_0.data}})[write_0.addr == 8'h55 & write_0_en];	// <stdin>:173:15, :939:12, :940:12, :941:12, :942:12, :943:12, :944:12, :946:12
  assign _T_169 = Register_inst85;	// <stdin>:946:12
  wire [31:0] _T_341 = ({{_T_168}, {write_0.data}})[write_0.addr == 8'h56 & write_0_en];	// <stdin>:172:15, :947:12, :948:12, :949:12, :950:12, :951:12, :952:12, :954:12
  assign _T_168 = Register_inst86;	// <stdin>:954:12
  wire [31:0] _T_342 = ({{_T_167}, {write_0.data}})[write_0.addr == 8'h57 & write_0_en];	// <stdin>:171:15, :955:12, :956:12, :957:12, :958:12, :959:12, :960:12, :962:12
  assign _T_167 = Register_inst87;	// <stdin>:962:12
  wire [31:0] _T_343 = ({{_T_166}, {write_0.data}})[write_0.addr == 8'h58 & write_0_en];	// <stdin>:170:15, :963:12, :964:12, :965:12, :966:12, :967:12, :968:12, :970:12
  assign _T_166 = Register_inst88;	// <stdin>:970:12
  wire [31:0] _T_344 = ({{_T_165}, {write_0.data}})[write_0.addr == 8'h59 & write_0_en];	// <stdin>:169:15, :971:12, :972:12, :973:12, :974:12, :975:12, :976:12, :978:12
  assign _T_165 = Register_inst89;	// <stdin>:978:12
  wire [31:0] _T_345 = ({{_T_164}, {write_0.data}})[write_0.addr == 8'h5A & write_0_en];	// <stdin>:168:15, :979:12, :980:12, :981:12, :982:12, :983:12, :984:12, :986:12
  assign _T_164 = Register_inst90;	// <stdin>:986:12
  wire [31:0] _T_346 = ({{_T_163}, {write_0.data}})[write_0.addr == 8'h5B & write_0_en];	// <stdin>:167:15, :987:12, :988:12, :989:12, :990:12, :991:12, :992:12, :994:12
  assign _T_163 = Register_inst91;	// <stdin>:994:12
  wire [31:0] _T_347 = ({{_T_162}, {write_0.data}})[write_0.addr == 8'h5C & write_0_en];	// <stdin>:166:15, :995:12, :996:12, :997:12, :998:12, :999:12, :1000:12, :1002:12
  assign _T_162 = Register_inst92;	// <stdin>:1002:12
  wire [31:0] _T_348 = ({{_T_161}, {write_0.data}})[write_0.addr == 8'h5D & write_0_en];	// <stdin>:165:15, :1003:12, :1004:12, :1005:12, :1006:12, :1007:12, :1008:12, :1010:12
  assign _T_161 = Register_inst93;	// <stdin>:1010:12
  wire [31:0] _T_349 = ({{_T_160}, {write_0.data}})[write_0.addr == 8'h5E & write_0_en];	// <stdin>:164:15, :1011:12, :1012:12, :1013:12, :1014:12, :1015:12, :1016:12, :1018:12
  assign _T_160 = Register_inst94;	// <stdin>:1018:12
  wire [31:0] _T_350 = ({{_T_159}, {write_0.data}})[write_0.addr == 8'h5F & write_0_en];	// <stdin>:163:15, :1019:12, :1020:12, :1021:12, :1022:12, :1023:12, :1024:12, :1026:12
  assign _T_159 = Register_inst95;	// <stdin>:1026:12
  wire [31:0] _T_351 = ({{_T_158}, {write_0.data}})[write_0.addr == 8'h60 & write_0_en];	// <stdin>:162:15, :1027:12, :1028:12, :1029:12, :1030:12, :1031:12, :1032:12, :1034:12
  assign _T_158 = Register_inst96;	// <stdin>:1034:12
  wire [31:0] _T_352 = ({{_T_157}, {write_0.data}})[write_0.addr == 8'h61 & write_0_en];	// <stdin>:161:15, :1035:12, :1036:12, :1037:12, :1038:12, :1039:12, :1040:12, :1042:12
  assign _T_157 = Register_inst97;	// <stdin>:1042:12
  wire [31:0] _T_353 = ({{_T_156}, {write_0.data}})[write_0.addr == 8'h62 & write_0_en];	// <stdin>:160:15, :1043:12, :1044:12, :1045:12, :1046:12, :1047:12, :1048:12, :1050:12
  assign _T_156 = Register_inst98;	// <stdin>:1050:12
  wire [31:0] _T_354 = ({{_T_155}, {write_0.data}})[write_0.addr == 8'h63 & write_0_en];	// <stdin>:159:15, :1051:12, :1052:12, :1053:12, :1054:12, :1055:12, :1056:12, :1058:12
  assign _T_155 = Register_inst99;	// <stdin>:1058:12
  wire [31:0] _T_355 = ({{_T_154}, {write_0.data}})[write_0.addr == 8'h64 & write_0_en];	// <stdin>:158:16, :1059:12, :1060:12, :1061:12, :1062:12, :1063:12, :1064:12, :1066:12
  assign _T_154 = Register_inst100;	// <stdin>:1066:12
  wire [31:0] _T_356 = ({{_T_153}, {write_0.data}})[write_0.addr == 8'h65 & write_0_en];	// <stdin>:157:16, :1067:12, :1068:12, :1069:12, :1070:12, :1071:12, :1072:12, :1074:12
  assign _T_153 = Register_inst101;	// <stdin>:1074:12
  wire [31:0] _T_357 = ({{_T_152}, {write_0.data}})[write_0.addr == 8'h66 & write_0_en];	// <stdin>:156:16, :1075:12, :1076:12, :1077:12, :1078:12, :1079:12, :1080:12, :1082:12
  assign _T_152 = Register_inst102;	// <stdin>:1082:12
  wire [31:0] _T_358 = ({{_T_151}, {write_0.data}})[write_0.addr == 8'h67 & write_0_en];	// <stdin>:155:16, :1083:12, :1084:12, :1085:12, :1086:12, :1087:12, :1088:12, :1090:12
  assign _T_151 = Register_inst103;	// <stdin>:1090:12
  wire [31:0] _T_359 = ({{_T_150}, {write_0.data}})[write_0.addr == 8'h68 & write_0_en];	// <stdin>:154:16, :1091:12, :1092:12, :1093:12, :1094:12, :1095:12, :1096:12, :1098:12
  assign _T_150 = Register_inst104;	// <stdin>:1098:12
  wire [31:0] _T_360 = ({{_T_149}, {write_0.data}})[write_0.addr == 8'h69 & write_0_en];	// <stdin>:153:16, :1099:12, :1100:12, :1101:12, :1102:12, :1103:12, :1104:12, :1106:12
  assign _T_149 = Register_inst105;	// <stdin>:1106:12
  wire [31:0] _T_361 = ({{_T_148}, {write_0.data}})[write_0.addr == 8'h6A & write_0_en];	// <stdin>:152:16, :1107:12, :1108:12, :1109:12, :1110:12, :1111:12, :1112:12, :1114:12
  assign _T_148 = Register_inst106;	// <stdin>:1114:12
  wire [31:0] _T_362 = ({{_T_147}, {write_0.data}})[write_0.addr == 8'h6B & write_0_en];	// <stdin>:151:16, :1115:12, :1116:12, :1117:12, :1118:12, :1119:12, :1120:12, :1122:12
  assign _T_147 = Register_inst107;	// <stdin>:1122:12
  wire [31:0] _T_363 = ({{_T_146}, {write_0.data}})[write_0.addr == 8'h6C & write_0_en];	// <stdin>:150:16, :1123:12, :1124:12, :1125:12, :1126:12, :1127:12, :1128:12, :1130:12
  assign _T_146 = Register_inst108;	// <stdin>:1130:12
  wire [31:0] _T_364 = ({{_T_145}, {write_0.data}})[write_0.addr == 8'h6D & write_0_en];	// <stdin>:149:16, :1131:12, :1132:12, :1133:12, :1134:12, :1135:12, :1136:12, :1138:12
  assign _T_145 = Register_inst109;	// <stdin>:1138:12
  wire [31:0] _T_365 = ({{_T_144}, {write_0.data}})[write_0.addr == 8'h6E & write_0_en];	// <stdin>:148:16, :1139:12, :1140:12, :1141:12, :1142:12, :1143:12, :1144:12, :1146:12
  assign _T_144 = Register_inst110;	// <stdin>:1146:12
  wire [31:0] _T_366 = ({{_T_143}, {write_0.data}})[write_0.addr == 8'h6F & write_0_en];	// <stdin>:147:16, :1147:12, :1148:12, :1149:12, :1150:12, :1151:12, :1152:12, :1154:12
  assign _T_143 = Register_inst111;	// <stdin>:1154:12
  wire [31:0] _T_367 = ({{_T_142}, {write_0.data}})[write_0.addr == 8'h70 & write_0_en];	// <stdin>:146:16, :1155:12, :1156:12, :1157:12, :1158:12, :1159:12, :1160:12, :1162:12
  assign _T_142 = Register_inst112;	// <stdin>:1162:12
  wire [31:0] _T_368 = ({{_T_141}, {write_0.data}})[write_0.addr == 8'h71 & write_0_en];	// <stdin>:145:16, :1163:12, :1164:12, :1165:12, :1166:12, :1167:12, :1168:12, :1170:12
  assign _T_141 = Register_inst113;	// <stdin>:1170:12
  wire [31:0] _T_369 = ({{_T_140}, {write_0.data}})[write_0.addr == 8'h72 & write_0_en];	// <stdin>:144:16, :1171:12, :1172:12, :1173:12, :1174:12, :1175:12, :1176:12, :1178:12
  assign _T_140 = Register_inst114;	// <stdin>:1178:12
  wire [31:0] _T_370 = ({{_T_139}, {write_0.data}})[write_0.addr == 8'h73 & write_0_en];	// <stdin>:143:16, :1179:12, :1180:12, :1181:12, :1182:12, :1183:12, :1184:12, :1186:12
  assign _T_139 = Register_inst115;	// <stdin>:1186:12
  wire [31:0] _T_371 = ({{_T_138}, {write_0.data}})[write_0.addr == 8'h74 & write_0_en];	// <stdin>:142:16, :1187:12, :1188:12, :1189:12, :1190:12, :1191:12, :1192:12, :1194:12
  assign _T_138 = Register_inst116;	// <stdin>:1194:12
  wire [31:0] _T_372 = ({{_T_137}, {write_0.data}})[write_0.addr == 8'h75 & write_0_en];	// <stdin>:141:16, :1195:12, :1196:12, :1197:12, :1198:12, :1199:12, :1200:12, :1202:12
  assign _T_137 = Register_inst117;	// <stdin>:1202:12
  wire [31:0] _T_373 = ({{_T_136}, {write_0.data}})[write_0.addr == 8'h76 & write_0_en];	// <stdin>:140:16, :1203:12, :1204:12, :1205:12, :1206:12, :1207:12, :1208:12, :1210:12
  assign _T_136 = Register_inst118;	// <stdin>:1210:12
  wire [31:0] _T_374 = ({{_T_135}, {write_0.data}})[write_0.addr == 8'h77 & write_0_en];	// <stdin>:139:16, :1211:12, :1212:12, :1213:12, :1214:12, :1215:12, :1216:12, :1218:12
  assign _T_135 = Register_inst119;	// <stdin>:1218:12
  wire [31:0] _T_375 = ({{_T_134}, {write_0.data}})[write_0.addr == 8'h78 & write_0_en];	// <stdin>:138:16, :1219:12, :1220:12, :1221:12, :1222:12, :1223:12, :1224:12, :1226:12
  assign _T_134 = Register_inst120;	// <stdin>:1226:12
  wire [31:0] _T_376 = ({{_T_133}, {write_0.data}})[write_0.addr == 8'h79 & write_0_en];	// <stdin>:137:16, :1227:12, :1228:12, :1229:12, :1230:12, :1231:12, :1232:12, :1234:12
  assign _T_133 = Register_inst121;	// <stdin>:1234:12
  wire [31:0] _T_377 = ({{_T_132}, {write_0.data}})[write_0.addr == 8'h7A & write_0_en];	// <stdin>:136:16, :1235:12, :1236:12, :1237:12, :1238:12, :1239:12, :1240:12, :1242:12
  assign _T_132 = Register_inst122;	// <stdin>:1242:12
  wire [31:0] _T_378 = ({{_T_131}, {write_0.data}})[write_0.addr == 8'h7B & write_0_en];	// <stdin>:135:16, :1243:12, :1244:12, :1245:12, :1246:12, :1247:12, :1248:12, :1250:12
  assign _T_131 = Register_inst123;	// <stdin>:1250:12
  wire [31:0] _T_379 = ({{_T_130}, {write_0.data}})[write_0.addr == 8'h7C & write_0_en];	// <stdin>:134:16, :1251:12, :1252:12, :1253:12, :1254:12, :1255:12, :1256:12, :1258:12
  assign _T_130 = Register_inst124;	// <stdin>:1258:12
  wire [31:0] _T_380 = ({{_T_129}, {write_0.data}})[write_0.addr == 8'h7D & write_0_en];	// <stdin>:133:16, :1259:12, :1260:12, :1261:12, :1262:12, :1263:12, :1264:12, :1266:12
  assign _T_129 = Register_inst125;	// <stdin>:1266:12
  wire [31:0] _T_381 = ({{_T_128}, {write_0.data}})[write_0.addr == 8'h7E & write_0_en];	// <stdin>:132:16, :1267:12, :1268:12, :1269:12, :1270:12, :1271:12, :1272:12, :1274:12
  assign _T_128 = Register_inst126;	// <stdin>:1274:12
  wire [31:0] _T_382 = ({{_T_127}, {write_0.data}})[write_0.addr == 8'h7F & write_0_en];	// <stdin>:131:16, :1275:12, :1276:12, :1277:12, :1278:12, :1279:12, :1280:12, :1282:12
  assign _T_127 = Register_inst127;	// <stdin>:1282:12
  wire [31:0] _T_383 = ({{_T_126}, {write_0.data}})[write_0.addr == 8'h80 & write_0_en];	// <stdin>:130:17, :1283:12, :1284:12, :1285:12, :1286:12, :1287:12, :1288:12, :1290:12
  assign _T_126 = Register_inst128;	// <stdin>:1290:12
  wire [31:0] _T_384 = ({{_T_125}, {write_0.data}})[write_0.addr == 8'h81 & write_0_en];	// <stdin>:129:17, :1291:12, :1292:12, :1293:12, :1294:12, :1295:12, :1296:12, :1298:12
  assign _T_125 = Register_inst129;	// <stdin>:1298:12
  wire [31:0] _T_385 = ({{_T_124}, {write_0.data}})[write_0.addr == 8'h82 & write_0_en];	// <stdin>:128:17, :1299:12, :1300:12, :1301:12, :1302:12, :1303:12, :1304:12, :1306:12
  assign _T_124 = Register_inst130;	// <stdin>:1306:12
  wire [31:0] _T_386 = ({{_T_123}, {write_0.data}})[write_0.addr == 8'h83 & write_0_en];	// <stdin>:127:17, :1307:12, :1308:12, :1309:12, :1310:12, :1311:12, :1312:12, :1314:12
  assign _T_123 = Register_inst131;	// <stdin>:1314:12
  wire [31:0] _T_387 = ({{_T_122}, {write_0.data}})[write_0.addr == 8'h84 & write_0_en];	// <stdin>:126:17, :1315:12, :1316:12, :1317:12, :1318:12, :1319:12, :1320:12, :1322:12
  assign _T_122 = Register_inst132;	// <stdin>:1322:12
  wire [31:0] _T_388 = ({{_T_121}, {write_0.data}})[write_0.addr == 8'h85 & write_0_en];	// <stdin>:125:17, :1323:12, :1324:12, :1325:12, :1326:12, :1327:12, :1328:12, :1330:12
  assign _T_121 = Register_inst133;	// <stdin>:1330:12
  wire [31:0] _T_389 = ({{_T_120}, {write_0.data}})[write_0.addr == 8'h86 & write_0_en];	// <stdin>:124:17, :1331:12, :1332:12, :1333:12, :1334:12, :1335:12, :1336:12, :1338:12
  assign _T_120 = Register_inst134;	// <stdin>:1338:12
  wire [31:0] _T_390 = ({{_T_119}, {write_0.data}})[write_0.addr == 8'h87 & write_0_en];	// <stdin>:123:17, :1339:12, :1340:12, :1341:12, :1342:12, :1343:12, :1344:12, :1346:12
  assign _T_119 = Register_inst135;	// <stdin>:1346:12
  wire [31:0] _T_391 = ({{_T_118}, {write_0.data}})[write_0.addr == 8'h88 & write_0_en];	// <stdin>:122:17, :1347:12, :1348:12, :1349:12, :1350:12, :1351:12, :1352:12, :1354:12
  assign _T_118 = Register_inst136;	// <stdin>:1354:12
  wire [31:0] _T_392 = ({{_T_117}, {write_0.data}})[write_0.addr == 8'h89 & write_0_en];	// <stdin>:121:17, :1355:12, :1356:12, :1357:12, :1358:12, :1359:12, :1360:12, :1362:12
  assign _T_117 = Register_inst137;	// <stdin>:1362:12
  wire [31:0] _T_393 = ({{_T_116}, {write_0.data}})[write_0.addr == 8'h8A & write_0_en];	// <stdin>:120:17, :1363:12, :1364:12, :1365:12, :1366:12, :1367:12, :1368:12, :1370:12
  assign _T_116 = Register_inst138;	// <stdin>:1370:12
  wire [31:0] _T_394 = ({{_T_115}, {write_0.data}})[write_0.addr == 8'h8B & write_0_en];	// <stdin>:119:17, :1371:12, :1372:12, :1373:12, :1374:12, :1375:12, :1376:12, :1378:12
  assign _T_115 = Register_inst139;	// <stdin>:1378:12
  wire [31:0] _T_395 = ({{_T_114}, {write_0.data}})[write_0.addr == 8'h8C & write_0_en];	// <stdin>:118:17, :1379:12, :1380:12, :1381:12, :1382:12, :1383:12, :1384:12, :1386:12
  assign _T_114 = Register_inst140;	// <stdin>:1386:12
  wire [31:0] _T_396 = ({{_T_113}, {write_0.data}})[write_0.addr == 8'h8D & write_0_en];	// <stdin>:117:17, :1387:12, :1388:12, :1389:12, :1390:12, :1391:12, :1392:12, :1394:12
  assign _T_113 = Register_inst141;	// <stdin>:1394:12
  wire [31:0] _T_397 = ({{_T_112}, {write_0.data}})[write_0.addr == 8'h8E & write_0_en];	// <stdin>:116:17, :1395:12, :1396:12, :1397:12, :1398:12, :1399:12, :1400:12, :1402:13
  assign _T_112 = Register_inst142;	// <stdin>:1402:13
  wire [31:0] _T_398 = ({{_T_111}, {write_0.data}})[write_0.addr == 8'h8F & write_0_en];	// <stdin>:115:17, :1403:13, :1404:13, :1405:13, :1406:13, :1407:13, :1408:13, :1410:13
  assign _T_111 = Register_inst143;	// <stdin>:1410:13
  wire [31:0] _T_399 = ({{_T_110}, {write_0.data}})[write_0.addr == 8'h90 & write_0_en];	// <stdin>:114:17, :1411:13, :1412:13, :1413:13, :1414:13, :1415:13, :1416:13, :1418:13
  assign _T_110 = Register_inst144;	// <stdin>:1418:13
  wire [31:0] _T_400 = ({{_T_109}, {write_0.data}})[write_0.addr == 8'h91 & write_0_en];	// <stdin>:113:17, :1419:13, :1420:13, :1421:13, :1422:13, :1423:13, :1424:13, :1426:13
  assign _T_109 = Register_inst145;	// <stdin>:1426:13
  wire [31:0] _T_401 = ({{_T_108}, {write_0.data}})[write_0.addr == 8'h92 & write_0_en];	// <stdin>:112:17, :1427:13, :1428:13, :1429:13, :1430:13, :1431:13, :1432:13, :1434:13
  assign _T_108 = Register_inst146;	// <stdin>:1434:13
  wire [31:0] _T_402 = ({{_T_107}, {write_0.data}})[write_0.addr == 8'h93 & write_0_en];	// <stdin>:111:17, :1435:13, :1436:13, :1437:13, :1438:13, :1439:13, :1440:13, :1442:13
  assign _T_107 = Register_inst147;	// <stdin>:1442:13
  wire [31:0] _T_403 = ({{_T_106}, {write_0.data}})[write_0.addr == 8'h94 & write_0_en];	// <stdin>:110:17, :1443:13, :1444:13, :1445:13, :1446:13, :1447:13, :1448:13, :1450:13
  assign _T_106 = Register_inst148;	// <stdin>:1450:13
  wire [31:0] _T_404 = ({{_T_105}, {write_0.data}})[write_0.addr == 8'h95 & write_0_en];	// <stdin>:109:17, :1451:13, :1452:13, :1453:13, :1454:13, :1455:13, :1456:13, :1458:13
  assign _T_105 = Register_inst149;	// <stdin>:1458:13
  wire [31:0] _T_405 = ({{_T_104}, {write_0.data}})[write_0.addr == 8'h96 & write_0_en];	// <stdin>:108:17, :1459:13, :1460:13, :1461:13, :1462:13, :1463:13, :1464:13, :1466:13
  assign _T_104 = Register_inst150;	// <stdin>:1466:13
  wire [31:0] _T_406 = ({{_T_103}, {write_0.data}})[write_0.addr == 8'h97 & write_0_en];	// <stdin>:107:17, :1467:13, :1468:13, :1469:13, :1470:13, :1471:13, :1472:13, :1474:13
  assign _T_103 = Register_inst151;	// <stdin>:1474:13
  wire [31:0] _T_407 = ({{_T_102}, {write_0.data}})[write_0.addr == 8'h98 & write_0_en];	// <stdin>:106:17, :1475:13, :1476:13, :1477:13, :1478:13, :1479:13, :1480:13, :1482:13
  assign _T_102 = Register_inst152;	// <stdin>:1482:13
  wire [31:0] _T_408 = ({{_T_101}, {write_0.data}})[write_0.addr == 8'h99 & write_0_en];	// <stdin>:105:17, :1483:13, :1484:13, :1485:13, :1486:13, :1487:13, :1488:13, :1490:13
  assign _T_101 = Register_inst153;	// <stdin>:1490:13
  wire [31:0] _T_409 = ({{_T_100}, {write_0.data}})[write_0.addr == 8'h9A & write_0_en];	// <stdin>:104:17, :1491:13, :1492:13, :1493:13, :1494:13, :1495:13, :1496:13, :1498:13
  assign _T_100 = Register_inst154;	// <stdin>:1498:13
  wire [31:0] _T_410 = ({{_T_99}, {write_0.data}})[write_0.addr == 8'h9B & write_0_en];	// <stdin>:103:17, :1499:13, :1500:13, :1501:13, :1502:13, :1503:13, :1504:13, :1506:13
  assign _T_99 = Register_inst155;	// <stdin>:1506:13
  wire [31:0] _T_411 = ({{_T_98}, {write_0.data}})[write_0.addr == 8'h9C & write_0_en];	// <stdin>:102:17, :1507:13, :1508:13, :1509:13, :1510:13, :1511:13, :1512:13, :1514:13
  assign _T_98 = Register_inst156;	// <stdin>:1514:13
  wire [31:0] _T_412 = ({{_T_97}, {write_0.data}})[write_0.addr == 8'h9D & write_0_en];	// <stdin>:101:16, :1515:13, :1516:13, :1517:13, :1518:13, :1519:13, :1520:13, :1522:13
  assign _T_97 = Register_inst157;	// <stdin>:1522:13
  wire [31:0] _T_413 = ({{_T_96}, {write_0.data}})[write_0.addr == 8'h9E & write_0_en];	// <stdin>:100:16, :1523:13, :1524:13, :1525:13, :1526:13, :1527:13, :1528:13, :1530:13
  assign _T_96 = Register_inst158;	// <stdin>:1530:13
  wire [31:0] _T_414 = ({{_T_95}, {write_0.data}})[write_0.addr == 8'h9F & write_0_en];	// <stdin>:99:16, :1531:13, :1532:13, :1533:13, :1534:13, :1535:13, :1536:13, :1538:13
  assign _T_95 = Register_inst159;	// <stdin>:1538:13
  wire [31:0] _T_415 = ({{_T_94}, {write_0.data}})[write_0.addr == 8'hA0 & write_0_en];	// <stdin>:98:16, :1539:13, :1540:13, :1541:13, :1542:13, :1543:13, :1544:13, :1546:13
  assign _T_94 = Register_inst160;	// <stdin>:1546:13
  wire [31:0] _T_416 = ({{_T_93}, {write_0.data}})[write_0.addr == 8'hA1 & write_0_en];	// <stdin>:97:16, :1547:13, :1548:13, :1549:13, :1550:13, :1551:13, :1552:13, :1554:13
  assign _T_93 = Register_inst161;	// <stdin>:1554:13
  wire [31:0] _T_417 = ({{_T_92}, {write_0.data}})[write_0.addr == 8'hA2 & write_0_en];	// <stdin>:96:16, :1555:13, :1556:13, :1557:13, :1558:13, :1559:13, :1560:13, :1562:13
  assign _T_92 = Register_inst162;	// <stdin>:1562:13
  wire [31:0] _T_418 = ({{_T_91}, {write_0.data}})[write_0.addr == 8'hA3 & write_0_en];	// <stdin>:95:16, :1563:13, :1564:13, :1565:13, :1566:13, :1567:13, :1568:13, :1570:13
  assign _T_91 = Register_inst163;	// <stdin>:1570:13
  wire [31:0] _T_419 = ({{_T_90}, {write_0.data}})[write_0.addr == 8'hA4 & write_0_en];	// <stdin>:94:16, :1571:13, :1572:13, :1573:13, :1574:13, :1575:13, :1576:13, :1578:13
  assign _T_90 = Register_inst164;	// <stdin>:1578:13
  wire [31:0] _T_420 = ({{_T_89}, {write_0.data}})[write_0.addr == 8'hA5 & write_0_en];	// <stdin>:93:16, :1579:13, :1580:13, :1581:13, :1582:13, :1583:13, :1584:13, :1586:13
  assign _T_89 = Register_inst165;	// <stdin>:1586:13
  wire [31:0] _T_421 = ({{_T_88}, {write_0.data}})[write_0.addr == 8'hA6 & write_0_en];	// <stdin>:92:16, :1587:13, :1588:13, :1589:13, :1590:13, :1591:13, :1592:13, :1594:13
  assign _T_88 = Register_inst166;	// <stdin>:1594:13
  wire [31:0] _T_422 = ({{_T_87}, {write_0.data}})[write_0.addr == 8'hA7 & write_0_en];	// <stdin>:91:16, :1595:13, :1596:13, :1597:13, :1598:13, :1599:13, :1600:13, :1602:13
  assign _T_87 = Register_inst167;	// <stdin>:1602:13
  wire [31:0] _T_423 = ({{_T_86}, {write_0.data}})[write_0.addr == 8'hA8 & write_0_en];	// <stdin>:90:16, :1603:13, :1604:13, :1605:13, :1606:13, :1607:13, :1608:13, :1610:13
  assign _T_86 = Register_inst168;	// <stdin>:1610:13
  wire [31:0] _T_424 = ({{_T_85}, {write_0.data}})[write_0.addr == 8'hA9 & write_0_en];	// <stdin>:89:16, :1611:13, :1612:13, :1613:13, :1614:13, :1615:13, :1616:13, :1618:13
  assign _T_85 = Register_inst169;	// <stdin>:1618:13
  wire [31:0] _T_425 = ({{_T_84}, {write_0.data}})[write_0.addr == 8'hAA & write_0_en];	// <stdin>:88:16, :1619:13, :1620:13, :1621:13, :1622:13, :1623:13, :1624:13, :1626:13
  assign _T_84 = Register_inst170;	// <stdin>:1626:13
  wire [31:0] _T_426 = ({{_T_83}, {write_0.data}})[write_0.addr == 8'hAB & write_0_en];	// <stdin>:87:16, :1627:13, :1628:13, :1629:13, :1630:13, :1631:13, :1632:13, :1634:13
  assign _T_83 = Register_inst171;	// <stdin>:1634:13
  wire [31:0] _T_427 = ({{_T_82}, {write_0.data}})[write_0.addr == 8'hAC & write_0_en];	// <stdin>:86:16, :1635:13, :1636:13, :1637:13, :1638:13, :1639:13, :1640:13, :1642:13
  assign _T_82 = Register_inst172;	// <stdin>:1642:13
  wire [31:0] _T_428 = ({{_T_81}, {write_0.data}})[write_0.addr == 8'hAD & write_0_en];	// <stdin>:85:16, :1643:13, :1644:13, :1645:13, :1646:13, :1647:13, :1648:13, :1650:13
  assign _T_81 = Register_inst173;	// <stdin>:1650:13
  wire [31:0] _T_429 = ({{_T_80}, {write_0.data}})[write_0.addr == 8'hAE & write_0_en];	// <stdin>:84:16, :1651:13, :1652:13, :1653:13, :1654:13, :1655:13, :1656:13, :1658:13
  assign _T_80 = Register_inst174;	// <stdin>:1658:13
  wire [31:0] _T_430 = ({{_T_79}, {write_0.data}})[write_0.addr == 8'hAF & write_0_en];	// <stdin>:83:16, :1659:13, :1660:13, :1661:13, :1662:13, :1663:13, :1664:13, :1666:13
  assign _T_79 = Register_inst175;	// <stdin>:1666:13
  wire [31:0] _T_431 = ({{_T_78}, {write_0.data}})[write_0.addr == 8'hB0 & write_0_en];	// <stdin>:82:16, :1667:13, :1668:13, :1669:13, :1670:13, :1671:13, :1672:13, :1674:13
  assign _T_78 = Register_inst176;	// <stdin>:1674:13
  wire [31:0] _T_432 = ({{_T_77}, {write_0.data}})[write_0.addr == 8'hB1 & write_0_en];	// <stdin>:81:16, :1675:13, :1676:13, :1677:13, :1678:13, :1679:13, :1680:13, :1682:13
  assign _T_77 = Register_inst177;	// <stdin>:1682:13
  wire [31:0] _T_433 = ({{_T_76}, {write_0.data}})[write_0.addr == 8'hB2 & write_0_en];	// <stdin>:80:16, :1683:13, :1684:13, :1685:13, :1686:13, :1687:13, :1688:13, :1690:13
  assign _T_76 = Register_inst178;	// <stdin>:1690:13
  wire [31:0] _T_434 = ({{_T_75}, {write_0.data}})[write_0.addr == 8'hB3 & write_0_en];	// <stdin>:79:16, :1691:13, :1692:13, :1693:13, :1694:13, :1695:13, :1696:13, :1698:13
  assign _T_75 = Register_inst179;	// <stdin>:1698:13
  wire [31:0] _T_435 = ({{_T_74}, {write_0.data}})[write_0.addr == 8'hB4 & write_0_en];	// <stdin>:78:16, :1699:13, :1700:13, :1701:13, :1702:13, :1703:13, :1704:13, :1706:13
  assign _T_74 = Register_inst180;	// <stdin>:1706:13
  wire [31:0] _T_436 = ({{_T_73}, {write_0.data}})[write_0.addr == 8'hB5 & write_0_en];	// <stdin>:77:16, :1707:13, :1708:13, :1709:13, :1710:13, :1711:13, :1712:13, :1714:13
  assign _T_73 = Register_inst181;	// <stdin>:1714:13
  wire [31:0] _T_437 = ({{_T_72}, {write_0.data}})[write_0.addr == 8'hB6 & write_0_en];	// <stdin>:76:16, :1715:13, :1716:13, :1717:13, :1718:13, :1719:13, :1720:13, :1722:13
  assign _T_72 = Register_inst182;	// <stdin>:1722:13
  wire [31:0] _T_438 = ({{_T_71}, {write_0.data}})[write_0.addr == 8'hB7 & write_0_en];	// <stdin>:75:16, :1723:13, :1724:13, :1725:13, :1726:13, :1727:13, :1728:13, :1730:13
  assign _T_71 = Register_inst183;	// <stdin>:1730:13
  wire [31:0] _T_439 = ({{_T_70}, {write_0.data}})[write_0.addr == 8'hB8 & write_0_en];	// <stdin>:74:16, :1731:13, :1732:13, :1733:13, :1734:13, :1735:13, :1736:13, :1738:13
  assign _T_70 = Register_inst184;	// <stdin>:1738:13
  wire [31:0] _T_440 = ({{_T_69}, {write_0.data}})[write_0.addr == 8'hB9 & write_0_en];	// <stdin>:73:16, :1739:13, :1740:13, :1741:13, :1742:13, :1743:13, :1744:13, :1746:13
  assign _T_69 = Register_inst185;	// <stdin>:1746:13
  wire [31:0] _T_441 = ({{_T_68}, {write_0.data}})[write_0.addr == 8'hBA & write_0_en];	// <stdin>:72:16, :1747:13, :1748:13, :1749:13, :1750:13, :1751:13, :1752:13, :1754:13
  assign _T_68 = Register_inst186;	// <stdin>:1754:13
  wire [31:0] _T_442 = ({{_T_67}, {write_0.data}})[write_0.addr == 8'hBB & write_0_en];	// <stdin>:71:16, :1755:13, :1756:13, :1757:13, :1758:13, :1759:13, :1760:13, :1762:13
  assign _T_67 = Register_inst187;	// <stdin>:1762:13
  wire [31:0] _T_443 = ({{_T_66}, {write_0.data}})[write_0.addr == 8'hBC & write_0_en];	// <stdin>:70:16, :1763:13, :1764:13, :1765:13, :1766:13, :1767:13, :1768:13, :1770:13
  assign _T_66 = Register_inst188;	// <stdin>:1770:13
  wire [31:0] _T_444 = ({{_T_65}, {write_0.data}})[write_0.addr == 8'hBD & write_0_en];	// <stdin>:69:16, :1771:13, :1772:13, :1773:13, :1774:13, :1775:13, :1776:13, :1778:13
  assign _T_65 = Register_inst189;	// <stdin>:1778:13
  wire [31:0] _T_445 = ({{_T_64}, {write_0.data}})[write_0.addr == 8'hBE & write_0_en];	// <stdin>:68:16, :1779:13, :1780:13, :1781:13, :1782:13, :1783:13, :1784:13, :1786:13
  assign _T_64 = Register_inst190;	// <stdin>:1786:13
  wire [31:0] _T_446 = ({{_T_63}, {write_0.data}})[write_0.addr == 8'hBF & write_0_en];	// <stdin>:67:16, :1787:13, :1788:13, :1789:13, :1790:13, :1791:13, :1792:13, :1794:13
  assign _T_63 = Register_inst191;	// <stdin>:1794:13
  wire [31:0] _T_447 = ({{_T_62}, {write_0.data}})[write_0.addr == 8'hC0 & write_0_en];	// <stdin>:66:16, :1795:13, :1796:13, :1797:13, :1798:13, :1799:13, :1800:13, :1802:13
  assign _T_62 = Register_inst192;	// <stdin>:1802:13
  wire [31:0] _T_448 = ({{_T_61}, {write_0.data}})[write_0.addr == 8'hC1 & write_0_en];	// <stdin>:65:16, :1803:13, :1804:13, :1805:13, :1806:13, :1807:13, :1808:13, :1810:13
  assign _T_61 = Register_inst193;	// <stdin>:1810:13
  wire [31:0] _T_449 = ({{_T_60}, {write_0.data}})[write_0.addr == 8'hC2 & write_0_en];	// <stdin>:64:16, :1811:13, :1812:13, :1813:13, :1814:13, :1815:13, :1816:13, :1818:13
  assign _T_60 = Register_inst194;	// <stdin>:1818:13
  wire [31:0] _T_450 = ({{_T_59}, {write_0.data}})[write_0.addr == 8'hC3 & write_0_en];	// <stdin>:63:16, :1819:13, :1820:13, :1821:13, :1822:13, :1823:13, :1824:13, :1826:13
  assign _T_59 = Register_inst195;	// <stdin>:1826:13
  wire [31:0] _T_451 = ({{_T_58}, {write_0.data}})[write_0.addr == 8'hC4 & write_0_en];	// <stdin>:62:16, :1827:13, :1828:13, :1829:13, :1830:13, :1831:13, :1832:13, :1834:13
  assign _T_58 = Register_inst196;	// <stdin>:1834:13
  wire [31:0] _T_452 = ({{_T_57}, {write_0.data}})[write_0.addr == 8'hC5 & write_0_en];	// <stdin>:61:16, :1835:13, :1836:13, :1837:13, :1838:13, :1839:13, :1840:13, :1842:13
  assign _T_57 = Register_inst197;	// <stdin>:1842:13
  wire [31:0] _T_453 = ({{_T_56}, {write_0.data}})[write_0.addr == 8'hC6 & write_0_en];	// <stdin>:60:16, :1843:13, :1844:13, :1845:13, :1846:13, :1847:13, :1848:13, :1850:13
  assign _T_56 = Register_inst198;	// <stdin>:1850:13
  wire [31:0] _T_454 = ({{_T_55}, {write_0.data}})[write_0.addr == 8'hC7 & write_0_en];	// <stdin>:59:16, :1851:13, :1852:13, :1853:13, :1854:13, :1855:13, :1856:13, :1858:13
  assign _T_55 = Register_inst199;	// <stdin>:1858:13
  wire [31:0] _T_455 = ({{_T_54}, {write_0.data}})[write_0.addr == 8'hC8 & write_0_en];	// <stdin>:58:16, :1859:13, :1860:13, :1861:13, :1862:13, :1863:13, :1864:13, :1866:13
  assign _T_54 = Register_inst200;	// <stdin>:1866:13
  wire [31:0] _T_456 = ({{_T_53}, {write_0.data}})[write_0.addr == 8'hC9 & write_0_en];	// <stdin>:57:16, :1867:13, :1868:13, :1869:13, :1870:13, :1871:13, :1872:13, :1874:13
  assign _T_53 = Register_inst201;	// <stdin>:1874:13
  wire [31:0] _T_457 = ({{_T_52}, {write_0.data}})[write_0.addr == 8'hCA & write_0_en];	// <stdin>:56:16, :1875:13, :1876:13, :1877:13, :1878:13, :1879:13, :1880:13, :1882:13
  assign _T_52 = Register_inst202;	// <stdin>:1882:13
  wire [31:0] _T_458 = ({{_T_51}, {write_0.data}})[write_0.addr == 8'hCB & write_0_en];	// <stdin>:55:16, :1883:13, :1884:13, :1885:13, :1886:13, :1887:13, :1888:13, :1890:13
  assign _T_51 = Register_inst203;	// <stdin>:1890:13
  wire [31:0] _T_459 = ({{_T_50}, {write_0.data}})[write_0.addr == 8'hCC & write_0_en];	// <stdin>:54:16, :1891:13, :1892:13, :1893:13, :1894:13, :1895:13, :1896:13, :1898:13
  assign _T_50 = Register_inst204;	// <stdin>:1898:13
  wire [31:0] _T_460 = ({{_T_49}, {write_0.data}})[write_0.addr == 8'hCD & write_0_en];	// <stdin>:53:16, :1899:13, :1900:13, :1901:13, :1902:13, :1903:13, :1904:13, :1906:13
  assign _T_49 = Register_inst205;	// <stdin>:1906:13
  wire [31:0] _T_461 = ({{_T_48}, {write_0.data}})[write_0.addr == 8'hCE & write_0_en];	// <stdin>:52:16, :1907:13, :1908:13, :1909:13, :1910:13, :1911:13, :1912:13, :1914:13
  assign _T_48 = Register_inst206;	// <stdin>:1914:13
  wire [31:0] _T_462 = ({{_T_47}, {write_0.data}})[write_0.addr == 8'hCF & write_0_en];	// <stdin>:51:16, :1915:13, :1916:13, :1917:13, :1918:13, :1919:13, :1920:13, :1922:13
  assign _T_47 = Register_inst207;	// <stdin>:1922:13
  wire [31:0] _T_463 = ({{_T_46}, {write_0.data}})[write_0.addr == 8'hD0 & write_0_en];	// <stdin>:50:16, :1923:13, :1924:13, :1925:13, :1926:13, :1927:13, :1928:13, :1930:13
  assign _T_46 = Register_inst208;	// <stdin>:1930:13
  wire [31:0] _T_464 = ({{_T_45}, {write_0.data}})[write_0.addr == 8'hD1 & write_0_en];	// <stdin>:49:16, :1931:13, :1932:13, :1933:13, :1934:13, :1935:13, :1936:13, :1938:13
  assign _T_45 = Register_inst209;	// <stdin>:1938:13
  wire [31:0] _T_465 = ({{_T_44}, {write_0.data}})[write_0.addr == 8'hD2 & write_0_en];	// <stdin>:48:16, :1939:13, :1940:13, :1941:13, :1942:13, :1943:13, :1944:13, :1946:13
  assign _T_44 = Register_inst210;	// <stdin>:1946:13
  wire [31:0] _T_466 = ({{_T_43}, {write_0.data}})[write_0.addr == 8'hD3 & write_0_en];	// <stdin>:47:16, :1947:13, :1948:13, :1949:13, :1950:13, :1951:13, :1952:13, :1954:13
  assign _T_43 = Register_inst211;	// <stdin>:1954:13
  wire [31:0] _T_467 = ({{_T_42}, {write_0.data}})[write_0.addr == 8'hD4 & write_0_en];	// <stdin>:46:16, :1955:13, :1956:13, :1957:13, :1958:13, :1959:13, :1960:13, :1962:13
  assign _T_42 = Register_inst212;	// <stdin>:1962:13
  wire [31:0] _T_468 = ({{_T_41}, {write_0.data}})[write_0.addr == 8'hD5 & write_0_en];	// <stdin>:45:16, :1963:13, :1964:13, :1965:13, :1966:13, :1967:13, :1968:13, :1970:13
  assign _T_41 = Register_inst213;	// <stdin>:1970:13
  wire [31:0] _T_469 = ({{_T_40}, {write_0.data}})[write_0.addr == 8'hD6 & write_0_en];	// <stdin>:44:16, :1971:13, :1972:13, :1973:13, :1974:13, :1975:13, :1976:13, :1978:13
  assign _T_40 = Register_inst214;	// <stdin>:1978:13
  wire [31:0] _T_470 = ({{_T_39}, {write_0.data}})[write_0.addr == 8'hD7 & write_0_en];	// <stdin>:43:16, :1979:13, :1980:13, :1981:13, :1982:13, :1983:13, :1984:13, :1986:13
  assign _T_39 = Register_inst215;	// <stdin>:1986:13
  wire [31:0] _T_471 = ({{_T_38}, {write_0.data}})[write_0.addr == 8'hD8 & write_0_en];	// <stdin>:42:16, :1987:13, :1988:13, :1989:13, :1990:13, :1991:13, :1992:13, :1994:13
  assign _T_38 = Register_inst216;	// <stdin>:1994:13
  wire [31:0] _T_472 = ({{_T_37}, {write_0.data}})[write_0.addr == 8'hD9 & write_0_en];	// <stdin>:41:16, :1995:13, :1996:13, :1997:13, :1998:13, :1999:13, :2000:13, :2002:13
  assign _T_37 = Register_inst217;	// <stdin>:2002:13
  wire [31:0] _T_473 = ({{_T_36}, {write_0.data}})[write_0.addr == 8'hDA & write_0_en];	// <stdin>:40:16, :2003:13, :2004:13, :2005:13, :2006:13, :2007:13, :2008:13, :2010:13
  assign _T_36 = Register_inst218;	// <stdin>:2010:13
  wire [31:0] _T_474 = ({{_T_35}, {write_0.data}})[write_0.addr == 8'hDB & write_0_en];	// <stdin>:39:16, :2011:13, :2012:13, :2013:13, :2014:13, :2015:13, :2016:13, :2018:13
  assign _T_35 = Register_inst219;	// <stdin>:2018:13
  wire [31:0] _T_475 = ({{_T_34}, {write_0.data}})[write_0.addr == 8'hDC & write_0_en];	// <stdin>:38:16, :2019:13, :2020:13, :2021:13, :2022:13, :2023:13, :2024:13, :2026:13
  assign _T_34 = Register_inst220;	// <stdin>:2026:13
  wire [31:0] _T_476 = ({{_T_33}, {write_0.data}})[write_0.addr == 8'hDD & write_0_en];	// <stdin>:37:16, :2027:13, :2028:13, :2029:13, :2030:13, :2031:13, :2032:13, :2034:13
  assign _T_33 = Register_inst221;	// <stdin>:2034:13
  wire [31:0] _T_477 = ({{_T_32}, {write_0.data}})[write_0.addr == 8'hDE & write_0_en];	// <stdin>:36:16, :2035:13, :2036:13, :2037:13, :2038:13, :2039:13, :2040:13, :2042:13
  assign _T_32 = Register_inst222;	// <stdin>:2042:13
  wire [31:0] _T_478 = ({{_T_31}, {write_0.data}})[write_0.addr == 8'hDF & write_0_en];	// <stdin>:35:16, :2043:13, :2044:13, :2045:13, :2046:13, :2047:13, :2048:13, :2050:13
  assign _T_31 = Register_inst223;	// <stdin>:2050:13
  wire [31:0] _T_479 = ({{_T_30}, {write_0.data}})[write_0.addr == 8'hE0 & write_0_en];	// <stdin>:34:16, :2051:13, :2052:13, :2053:13, :2054:13, :2055:13, :2056:13, :2058:13
  assign _T_30 = Register_inst224;	// <stdin>:2058:13
  wire [31:0] _T_480 = ({{_T_29}, {write_0.data}})[write_0.addr == 8'hE1 & write_0_en];	// <stdin>:33:16, :2059:13, :2060:13, :2061:13, :2062:13, :2063:13, :2064:13, :2066:13
  assign _T_29 = Register_inst225;	// <stdin>:2066:13
  wire [31:0] _T_481 = ({{_T_28}, {write_0.data}})[write_0.addr == 8'hE2 & write_0_en];	// <stdin>:32:16, :2067:13, :2068:13, :2069:13, :2070:13, :2071:13, :2072:13, :2074:13
  assign _T_28 = Register_inst226;	// <stdin>:2074:13
  wire [31:0] _T_482 = ({{_T_27}, {write_0.data}})[write_0.addr == 8'hE3 & write_0_en];	// <stdin>:31:16, :2075:13, :2076:13, :2077:13, :2078:13, :2079:13, :2080:13, :2082:13
  assign _T_27 = Register_inst227;	// <stdin>:2082:13
  wire [31:0] _T_483 = ({{_T_26}, {write_0.data}})[write_0.addr == 8'hE4 & write_0_en];	// <stdin>:30:16, :2083:13, :2084:13, :2085:13, :2086:13, :2087:13, :2088:13, :2090:13
  assign _T_26 = Register_inst228;	// <stdin>:2090:13
  wire [31:0] _T_484 = ({{_T_25}, {write_0.data}})[write_0.addr == 8'hE5 & write_0_en];	// <stdin>:29:16, :2091:13, :2092:13, :2093:13, :2094:13, :2095:13, :2096:13, :2098:13
  assign _T_25 = Register_inst229;	// <stdin>:2098:13
  wire [31:0] _T_485 = ({{_T_24}, {write_0.data}})[write_0.addr == 8'hE6 & write_0_en];	// <stdin>:28:16, :2099:13, :2100:13, :2101:13, :2102:13, :2103:13, :2104:13, :2106:13
  assign _T_24 = Register_inst230;	// <stdin>:2106:13
  wire [31:0] _T_486 = ({{_T_23}, {write_0.data}})[write_0.addr == 8'hE7 & write_0_en];	// <stdin>:27:16, :2107:13, :2108:13, :2109:13, :2110:13, :2111:13, :2112:13, :2114:13
  assign _T_23 = Register_inst231;	// <stdin>:2114:13
  wire [31:0] _T_487 = ({{_T_22}, {write_0.data}})[write_0.addr == 8'hE8 & write_0_en];	// <stdin>:26:16, :2115:13, :2116:13, :2117:13, :2118:13, :2119:13, :2120:13, :2122:13
  assign _T_22 = Register_inst232;	// <stdin>:2122:13
  wire [31:0] _T_488 = ({{_T_21}, {write_0.data}})[write_0.addr == 8'hE9 & write_0_en];	// <stdin>:25:16, :2123:13, :2124:13, :2125:13, :2126:13, :2127:13, :2128:13, :2130:13
  assign _T_21 = Register_inst233;	// <stdin>:2130:13
  wire [31:0] _T_489 = ({{_T_20}, {write_0.data}})[write_0.addr == 8'hEA & write_0_en];	// <stdin>:24:16, :2131:13, :2132:13, :2133:13, :2134:13, :2135:13, :2136:13, :2138:13
  assign _T_20 = Register_inst234;	// <stdin>:2138:13
  wire [31:0] _T_490 = ({{_T_19}, {write_0.data}})[write_0.addr == 8'hEB & write_0_en];	// <stdin>:23:16, :2139:13, :2140:13, :2141:13, :2142:13, :2143:13, :2144:13, :2146:13
  assign _T_19 = Register_inst235;	// <stdin>:2146:13
  wire [31:0] _T_491 = ({{_T_18}, {write_0.data}})[write_0.addr == 8'hEC & write_0_en];	// <stdin>:22:16, :2147:13, :2148:13, :2149:13, :2150:13, :2151:13, :2152:13, :2154:13
  assign _T_18 = Register_inst236;	// <stdin>:2154:13
  wire [31:0] _T_492 = ({{_T_17}, {write_0.data}})[write_0.addr == 8'hED & write_0_en];	// <stdin>:21:16, :2155:13, :2156:13, :2157:13, :2158:13, :2159:13, :2160:13, :2162:13
  assign _T_17 = Register_inst237;	// <stdin>:2162:13
  wire [31:0] _T_493 = ({{_T_16}, {write_0.data}})[write_0.addr == 8'hEE & write_0_en];	// <stdin>:20:16, :2163:13, :2164:13, :2165:13, :2166:13, :2167:13, :2168:13, :2170:13
  assign _T_16 = Register_inst238;	// <stdin>:2170:13
  wire [31:0] _T_494 = ({{_T_15}, {write_0.data}})[write_0.addr == 8'hEF & write_0_en];	// <stdin>:19:16, :2171:13, :2172:13, :2173:13, :2174:13, :2175:13, :2176:13, :2178:13
  assign _T_15 = Register_inst239;	// <stdin>:2178:13
  wire [31:0] _T_495 = ({{_T_14}, {write_0.data}})[write_0.addr == 8'hF0 & write_0_en];	// <stdin>:18:16, :2179:13, :2180:13, :2181:13, :2182:13, :2183:13, :2184:13, :2186:13
  assign _T_14 = Register_inst240;	// <stdin>:2186:13
  wire [31:0] _T_496 = ({{_T_13}, {write_0.data}})[write_0.addr == 8'hF1 & write_0_en];	// <stdin>:17:16, :2187:13, :2188:13, :2189:13, :2190:13, :2191:13, :2192:13, :2194:13
  assign _T_13 = Register_inst241;	// <stdin>:2194:13
  wire [31:0] _T_497 = ({{_T_12}, {write_0.data}})[write_0.addr == 8'hF2 & write_0_en];	// <stdin>:16:16, :2195:13, :2196:13, :2197:13, :2198:13, :2199:13, :2200:13, :2202:13
  assign _T_12 = Register_inst242;	// <stdin>:2202:13
  wire [31:0] _T_498 = ({{_T_11}, {write_0.data}})[write_0.addr == 8'hF3 & write_0_en];	// <stdin>:15:16, :2203:13, :2204:13, :2205:13, :2206:13, :2207:13, :2208:13, :2210:13
  assign _T_11 = Register_inst243;	// <stdin>:2210:13
  wire [31:0] _T_499 = ({{_T_10}, {write_0.data}})[write_0.addr == 8'hF4 & write_0_en];	// <stdin>:14:16, :2211:13, :2212:13, :2213:13, :2214:13, :2215:13, :2216:13, :2218:13
  assign _T_10 = Register_inst244;	// <stdin>:2218:13
  wire [31:0] _T_500 = ({{_T_9}, {write_0.data}})[write_0.addr == 8'hF5 & write_0_en];	// <stdin>:13:16, :2219:13, :2220:13, :2221:13, :2222:13, :2223:13, :2224:13, :2226:13
  assign _T_9 = Register_inst245;	// <stdin>:2226:13
  wire [31:0] _T_501 = ({{_T_8}, {write_0.data}})[write_0.addr == 8'hF6 & write_0_en];	// <stdin>:12:16, :2227:13, :2228:13, :2229:13, :2230:13, :2231:13, :2232:13, :2234:13
  assign _T_8 = Register_inst246;	// <stdin>:2234:13
  wire [31:0] _T_502 = ({{_T_7}, {write_0.data}})[write_0.addr == 8'hF7 & write_0_en];	// <stdin>:11:15, :2235:13, :2236:13, :2237:13, :2238:13, :2239:13, :2240:13, :2242:13
  assign _T_7 = Register_inst247;	// <stdin>:2242:13
  wire [31:0] _T_503 = ({{_T_6}, {write_0.data}})[write_0.addr == 8'hF8 & write_0_en];	// <stdin>:10:15, :2243:13, :2244:13, :2245:13, :2246:13, :2247:13, :2248:13, :2250:13
  assign _T_6 = Register_inst248;	// <stdin>:2250:13
  wire [31:0] _T_504 = ({{_T_5}, {write_0.data}})[write_0.addr == 8'hF9 & write_0_en];	// <stdin>:9:15, :2251:13, :2252:13, :2253:13, :2254:13, :2255:13, :2256:13, :2258:13
  assign _T_5 = Register_inst249;	// <stdin>:2258:13
  wire [31:0] _T_505 = ({{_T_4}, {write_0.data}})[write_0.addr == 8'hFA & write_0_en];	// <stdin>:8:15, :2259:13, :2260:13, :2261:13, :2262:13, :2263:13, :2264:13, :2266:13
  assign _T_4 = Register_inst250;	// <stdin>:2266:13
  wire [31:0] _T_506 = ({{_T_3}, {write_0.data}})[write_0.addr == 8'hFB & write_0_en];	// <stdin>:7:15, :2267:13, :2268:13, :2269:13, :2270:13, :2271:13, :2272:13, :2274:13
  assign _T_3 = Register_inst251;	// <stdin>:2274:13
  wire [31:0] _T_507 = ({{_T_2}, {write_0.data}})[write_0.addr == 8'hFC & write_0_en];	// <stdin>:6:15, :2275:13, :2276:13, :2277:13, :2278:13, :2279:13, :2280:13, :2282:13
  assign _T_2 = Register_inst252;	// <stdin>:2282:13
  wire [31:0] _T_508 = ({{_T_1}, {write_0.data}})[write_0.addr == 8'hFD & write_0_en];	// <stdin>:5:15, :2283:13, :2284:13, :2285:13, :2286:13, :2287:13, :2288:13, :2290:13
  assign _T_1 = Register_inst253;	// <stdin>:2290:13
  wire [31:0] _T_509 = ({{_T_0}, {write_0.data}})[write_0.addr == 8'hFE & write_0_en];	// <stdin>:4:15, :2291:13, :2292:13, :2293:13, :2294:13, :2295:13, :2296:13, :2298:13
  assign _T_0 = Register_inst254;	// <stdin>:2298:13
  wire [31:0] _T_510 = ({{_T}, {write_0.data}})[&write_0.addr & write_0_en];	// <stdin>:2299:13, :2300:13, :2301:13, :2302:13, :2303:13, :2304:13, :3081:13
  always @(posedge CLK or posedge ASYNCRESET) begin	// <stdin>:2306:5
    if (ASYNCRESET) begin	// <stdin>:2306:5
      Register_inst0 <= 32'h0;	// <stdin>:2564:17, :2565:7
      Register_inst1 <= 32'h0;	// <stdin>:2564:17, :2566:7
      Register_inst2 <= 32'h0;	// <stdin>:2564:17, :2567:7
      Register_inst3 <= 32'h0;	// <stdin>:2564:17, :2568:7
      Register_inst4 <= 32'h0;	// <stdin>:2564:17, :2569:7
      Register_inst5 <= 32'h0;	// <stdin>:2564:17, :2570:7
      Register_inst6 <= 32'h0;	// <stdin>:2564:17, :2571:7
      Register_inst7 <= 32'h0;	// <stdin>:2564:17, :2572:7
      Register_inst8 <= 32'h0;	// <stdin>:2564:17, :2573:7
      Register_inst9 <= 32'h0;	// <stdin>:2564:17, :2574:7
      Register_inst10 <= 32'h0;	// <stdin>:2564:17, :2575:7
      Register_inst11 <= 32'h0;	// <stdin>:2564:17, :2576:7
      Register_inst12 <= 32'h0;	// <stdin>:2564:17, :2577:7
      Register_inst13 <= 32'h0;	// <stdin>:2564:17, :2578:7
      Register_inst14 <= 32'h0;	// <stdin>:2564:17, :2579:7
      Register_inst15 <= 32'h0;	// <stdin>:2564:17, :2580:7
      Register_inst16 <= 32'h0;	// <stdin>:2564:17, :2581:7
      Register_inst17 <= 32'h0;	// <stdin>:2564:17, :2582:7
      Register_inst18 <= 32'h0;	// <stdin>:2564:17, :2583:7
      Register_inst19 <= 32'h0;	// <stdin>:2564:17, :2584:7
      Register_inst20 <= 32'h0;	// <stdin>:2564:17, :2585:7
      Register_inst21 <= 32'h0;	// <stdin>:2564:17, :2586:7
      Register_inst22 <= 32'h0;	// <stdin>:2564:17, :2587:7
      Register_inst23 <= 32'h0;	// <stdin>:2564:17, :2588:7
      Register_inst24 <= 32'h0;	// <stdin>:2564:17, :2589:7
      Register_inst25 <= 32'h0;	// <stdin>:2564:17, :2590:7
      Register_inst26 <= 32'h0;	// <stdin>:2564:17, :2591:7
      Register_inst27 <= 32'h0;	// <stdin>:2564:17, :2592:7
      Register_inst28 <= 32'h0;	// <stdin>:2564:17, :2593:7
      Register_inst29 <= 32'h0;	// <stdin>:2564:17, :2594:7
      Register_inst30 <= 32'h0;	// <stdin>:2564:17, :2595:7
      Register_inst31 <= 32'h0;	// <stdin>:2564:17, :2596:7
      Register_inst32 <= 32'h0;	// <stdin>:2564:17, :2597:7
      Register_inst33 <= 32'h0;	// <stdin>:2564:17, :2598:7
      Register_inst34 <= 32'h0;	// <stdin>:2564:17, :2599:7
      Register_inst35 <= 32'h0;	// <stdin>:2564:17, :2600:7
      Register_inst36 <= 32'h0;	// <stdin>:2564:17, :2601:7
      Register_inst37 <= 32'h0;	// <stdin>:2564:17, :2602:7
      Register_inst38 <= 32'h0;	// <stdin>:2564:17, :2603:7
      Register_inst39 <= 32'h0;	// <stdin>:2564:17, :2604:7
      Register_inst40 <= 32'h0;	// <stdin>:2564:17, :2605:7
      Register_inst41 <= 32'h0;	// <stdin>:2564:17, :2606:7
      Register_inst42 <= 32'h0;	// <stdin>:2564:17, :2607:7
      Register_inst43 <= 32'h0;	// <stdin>:2564:17, :2608:7
      Register_inst44 <= 32'h0;	// <stdin>:2564:17, :2609:7
      Register_inst45 <= 32'h0;	// <stdin>:2564:17, :2610:7
      Register_inst46 <= 32'h0;	// <stdin>:2564:17, :2611:7
      Register_inst47 <= 32'h0;	// <stdin>:2564:17, :2612:7
      Register_inst48 <= 32'h0;	// <stdin>:2564:17, :2613:7
      Register_inst49 <= 32'h0;	// <stdin>:2564:17, :2614:7
      Register_inst50 <= 32'h0;	// <stdin>:2564:17, :2615:7
      Register_inst51 <= 32'h0;	// <stdin>:2564:17, :2616:7
      Register_inst52 <= 32'h0;	// <stdin>:2564:17, :2617:7
      Register_inst53 <= 32'h0;	// <stdin>:2564:17, :2618:7
      Register_inst54 <= 32'h0;	// <stdin>:2564:17, :2619:7
      Register_inst55 <= 32'h0;	// <stdin>:2564:17, :2620:7
      Register_inst56 <= 32'h0;	// <stdin>:2564:17, :2621:7
      Register_inst57 <= 32'h0;	// <stdin>:2564:17, :2622:7
      Register_inst58 <= 32'h0;	// <stdin>:2564:17, :2623:7
      Register_inst59 <= 32'h0;	// <stdin>:2564:17, :2624:7
      Register_inst60 <= 32'h0;	// <stdin>:2564:17, :2625:7
      Register_inst61 <= 32'h0;	// <stdin>:2564:17, :2626:7
      Register_inst62 <= 32'h0;	// <stdin>:2564:17, :2627:7
      Register_inst63 <= 32'h0;	// <stdin>:2564:17, :2628:7
      Register_inst64 <= 32'h0;	// <stdin>:2564:17, :2629:7
      Register_inst65 <= 32'h0;	// <stdin>:2564:17, :2630:7
      Register_inst66 <= 32'h0;	// <stdin>:2564:17, :2631:7
      Register_inst67 <= 32'h0;	// <stdin>:2564:17, :2632:7
      Register_inst68 <= 32'h0;	// <stdin>:2564:17, :2633:7
      Register_inst69 <= 32'h0;	// <stdin>:2564:17, :2634:7
      Register_inst70 <= 32'h0;	// <stdin>:2564:17, :2635:7
      Register_inst71 <= 32'h0;	// <stdin>:2564:17, :2636:7
      Register_inst72 <= 32'h0;	// <stdin>:2564:17, :2637:7
      Register_inst73 <= 32'h0;	// <stdin>:2564:17, :2638:7
      Register_inst74 <= 32'h0;	// <stdin>:2564:17, :2639:7
      Register_inst75 <= 32'h0;	// <stdin>:2564:17, :2640:7
      Register_inst76 <= 32'h0;	// <stdin>:2564:17, :2641:7
      Register_inst77 <= 32'h0;	// <stdin>:2564:17, :2642:7
      Register_inst78 <= 32'h0;	// <stdin>:2564:17, :2643:7
      Register_inst79 <= 32'h0;	// <stdin>:2564:17, :2644:7
      Register_inst80 <= 32'h0;	// <stdin>:2564:17, :2645:7
      Register_inst81 <= 32'h0;	// <stdin>:2564:17, :2646:7
      Register_inst82 <= 32'h0;	// <stdin>:2564:17, :2647:7
      Register_inst83 <= 32'h0;	// <stdin>:2564:17, :2648:7
      Register_inst84 <= 32'h0;	// <stdin>:2564:17, :2649:7
      Register_inst85 <= 32'h0;	// <stdin>:2564:17, :2650:7
      Register_inst86 <= 32'h0;	// <stdin>:2564:17, :2651:7
      Register_inst87 <= 32'h0;	// <stdin>:2564:17, :2652:7
      Register_inst88 <= 32'h0;	// <stdin>:2564:17, :2653:7
      Register_inst89 <= 32'h0;	// <stdin>:2564:17, :2654:7
      Register_inst90 <= 32'h0;	// <stdin>:2564:17, :2655:7
      Register_inst91 <= 32'h0;	// <stdin>:2564:17, :2656:7
      Register_inst92 <= 32'h0;	// <stdin>:2564:17, :2657:7
      Register_inst93 <= 32'h0;	// <stdin>:2564:17, :2658:7
      Register_inst94 <= 32'h0;	// <stdin>:2564:17, :2659:7
      Register_inst95 <= 32'h0;	// <stdin>:2564:17, :2660:7
      Register_inst96 <= 32'h0;	// <stdin>:2564:17, :2661:7
      Register_inst97 <= 32'h0;	// <stdin>:2564:17, :2662:7
      Register_inst98 <= 32'h0;	// <stdin>:2564:17, :2663:7
      Register_inst99 <= 32'h0;	// <stdin>:2564:17, :2664:7
      Register_inst100 <= 32'h0;	// <stdin>:2564:17, :2665:7
      Register_inst101 <= 32'h0;	// <stdin>:2564:17, :2666:7
      Register_inst102 <= 32'h0;	// <stdin>:2564:17, :2667:7
      Register_inst103 <= 32'h0;	// <stdin>:2564:17, :2668:7
      Register_inst104 <= 32'h0;	// <stdin>:2564:17, :2669:7
      Register_inst105 <= 32'h0;	// <stdin>:2564:17, :2670:7
      Register_inst106 <= 32'h0;	// <stdin>:2564:17, :2671:7
      Register_inst107 <= 32'h0;	// <stdin>:2564:17, :2672:7
      Register_inst108 <= 32'h0;	// <stdin>:2564:17, :2673:7
      Register_inst109 <= 32'h0;	// <stdin>:2564:17, :2674:7
      Register_inst110 <= 32'h0;	// <stdin>:2564:17, :2675:7
      Register_inst111 <= 32'h0;	// <stdin>:2564:17, :2676:7
      Register_inst112 <= 32'h0;	// <stdin>:2564:17, :2677:7
      Register_inst113 <= 32'h0;	// <stdin>:2564:17, :2678:7
      Register_inst114 <= 32'h0;	// <stdin>:2564:17, :2679:7
      Register_inst115 <= 32'h0;	// <stdin>:2564:17, :2680:7
      Register_inst116 <= 32'h0;	// <stdin>:2564:17, :2681:7
      Register_inst117 <= 32'h0;	// <stdin>:2564:17, :2682:7
      Register_inst118 <= 32'h0;	// <stdin>:2564:17, :2683:7
      Register_inst119 <= 32'h0;	// <stdin>:2564:17, :2684:7
      Register_inst120 <= 32'h0;	// <stdin>:2564:17, :2685:7
      Register_inst121 <= 32'h0;	// <stdin>:2564:17, :2686:7
      Register_inst122 <= 32'h0;	// <stdin>:2564:17, :2687:7
      Register_inst123 <= 32'h0;	// <stdin>:2564:17, :2688:7
      Register_inst124 <= 32'h0;	// <stdin>:2564:17, :2689:7
      Register_inst125 <= 32'h0;	// <stdin>:2564:17, :2690:7
      Register_inst126 <= 32'h0;	// <stdin>:2564:17, :2691:7
      Register_inst127 <= 32'h0;	// <stdin>:2564:17, :2692:7
      Register_inst128 <= 32'h0;	// <stdin>:2564:17, :2693:7
      Register_inst129 <= 32'h0;	// <stdin>:2564:17, :2694:7
      Register_inst130 <= 32'h0;	// <stdin>:2564:17, :2695:7
      Register_inst131 <= 32'h0;	// <stdin>:2564:17, :2696:7
      Register_inst132 <= 32'h0;	// <stdin>:2564:17, :2697:7
      Register_inst133 <= 32'h0;	// <stdin>:2564:17, :2698:7
      Register_inst134 <= 32'h0;	// <stdin>:2564:17, :2699:7
      Register_inst135 <= 32'h0;	// <stdin>:2564:17, :2700:7
      Register_inst136 <= 32'h0;	// <stdin>:2564:17, :2701:7
      Register_inst137 <= 32'h0;	// <stdin>:2564:17, :2702:7
      Register_inst138 <= 32'h0;	// <stdin>:2564:17, :2703:7
      Register_inst139 <= 32'h0;	// <stdin>:2564:17, :2704:7
      Register_inst140 <= 32'h0;	// <stdin>:2564:17, :2705:7
      Register_inst141 <= 32'h0;	// <stdin>:2564:17, :2706:7
      Register_inst142 <= 32'h0;	// <stdin>:2564:17, :2707:7
      Register_inst143 <= 32'h0;	// <stdin>:2564:17, :2708:7
      Register_inst144 <= 32'h0;	// <stdin>:2564:17, :2709:7
      Register_inst145 <= 32'h0;	// <stdin>:2564:17, :2710:7
      Register_inst146 <= 32'h0;	// <stdin>:2564:17, :2711:7
      Register_inst147 <= 32'h0;	// <stdin>:2564:17, :2712:7
      Register_inst148 <= 32'h0;	// <stdin>:2564:17, :2713:7
      Register_inst149 <= 32'h0;	// <stdin>:2564:17, :2714:7
      Register_inst150 <= 32'h0;	// <stdin>:2564:17, :2715:7
      Register_inst151 <= 32'h0;	// <stdin>:2564:17, :2716:7
      Register_inst152 <= 32'h0;	// <stdin>:2564:17, :2717:7
      Register_inst153 <= 32'h0;	// <stdin>:2564:17, :2718:7
      Register_inst154 <= 32'h0;	// <stdin>:2564:17, :2719:7
      Register_inst155 <= 32'h0;	// <stdin>:2564:17, :2720:7
      Register_inst156 <= 32'h0;	// <stdin>:2564:17, :2721:7
      Register_inst157 <= 32'h0;	// <stdin>:2564:17, :2722:7
      Register_inst158 <= 32'h0;	// <stdin>:2564:17, :2723:7
      Register_inst159 <= 32'h0;	// <stdin>:2564:17, :2724:7
      Register_inst160 <= 32'h0;	// <stdin>:2564:17, :2725:7
      Register_inst161 <= 32'h0;	// <stdin>:2564:17, :2726:7
      Register_inst162 <= 32'h0;	// <stdin>:2564:17, :2727:7
      Register_inst163 <= 32'h0;	// <stdin>:2564:17, :2728:7
      Register_inst164 <= 32'h0;	// <stdin>:2564:17, :2729:7
      Register_inst165 <= 32'h0;	// <stdin>:2564:17, :2730:7
      Register_inst166 <= 32'h0;	// <stdin>:2564:17, :2731:7
      Register_inst167 <= 32'h0;	// <stdin>:2564:17, :2732:7
      Register_inst168 <= 32'h0;	// <stdin>:2564:17, :2733:7
      Register_inst169 <= 32'h0;	// <stdin>:2564:17, :2734:7
      Register_inst170 <= 32'h0;	// <stdin>:2564:17, :2735:7
      Register_inst171 <= 32'h0;	// <stdin>:2564:17, :2736:7
      Register_inst172 <= 32'h0;	// <stdin>:2564:17, :2737:7
      Register_inst173 <= 32'h0;	// <stdin>:2564:17, :2738:7
      Register_inst174 <= 32'h0;	// <stdin>:2564:17, :2739:7
      Register_inst175 <= 32'h0;	// <stdin>:2564:17, :2740:7
      Register_inst176 <= 32'h0;	// <stdin>:2564:17, :2741:7
      Register_inst177 <= 32'h0;	// <stdin>:2564:17, :2742:7
      Register_inst178 <= 32'h0;	// <stdin>:2564:17, :2743:7
      Register_inst179 <= 32'h0;	// <stdin>:2564:17, :2744:7
      Register_inst180 <= 32'h0;	// <stdin>:2564:17, :2745:7
      Register_inst181 <= 32'h0;	// <stdin>:2564:17, :2746:7
      Register_inst182 <= 32'h0;	// <stdin>:2564:17, :2747:7
      Register_inst183 <= 32'h0;	// <stdin>:2564:17, :2748:7
      Register_inst184 <= 32'h0;	// <stdin>:2564:17, :2749:7
      Register_inst185 <= 32'h0;	// <stdin>:2564:17, :2750:7
      Register_inst186 <= 32'h0;	// <stdin>:2564:17, :2751:7
      Register_inst187 <= 32'h0;	// <stdin>:2564:17, :2752:7
      Register_inst188 <= 32'h0;	// <stdin>:2564:17, :2753:7
      Register_inst189 <= 32'h0;	// <stdin>:2564:17, :2754:7
      Register_inst190 <= 32'h0;	// <stdin>:2564:17, :2755:7
      Register_inst191 <= 32'h0;	// <stdin>:2564:17, :2756:7
      Register_inst192 <= 32'h0;	// <stdin>:2564:17, :2757:7
      Register_inst193 <= 32'h0;	// <stdin>:2564:17, :2758:7
      Register_inst194 <= 32'h0;	// <stdin>:2564:17, :2759:7
      Register_inst195 <= 32'h0;	// <stdin>:2564:17, :2760:7
      Register_inst196 <= 32'h0;	// <stdin>:2564:17, :2761:7
      Register_inst197 <= 32'h0;	// <stdin>:2564:17, :2762:7
      Register_inst198 <= 32'h0;	// <stdin>:2564:17, :2763:7
      Register_inst199 <= 32'h0;	// <stdin>:2564:17, :2764:7
      Register_inst200 <= 32'h0;	// <stdin>:2564:17, :2765:7
      Register_inst201 <= 32'h0;	// <stdin>:2564:17, :2766:7
      Register_inst202 <= 32'h0;	// <stdin>:2564:17, :2767:7
      Register_inst203 <= 32'h0;	// <stdin>:2564:17, :2768:7
      Register_inst204 <= 32'h0;	// <stdin>:2564:17, :2769:7
      Register_inst205 <= 32'h0;	// <stdin>:2564:17, :2770:7
      Register_inst206 <= 32'h0;	// <stdin>:2564:17, :2771:7
      Register_inst207 <= 32'h0;	// <stdin>:2564:17, :2772:7
      Register_inst208 <= 32'h0;	// <stdin>:2564:17, :2773:7
      Register_inst209 <= 32'h0;	// <stdin>:2564:17, :2774:7
      Register_inst210 <= 32'h0;	// <stdin>:2564:17, :2775:7
      Register_inst211 <= 32'h0;	// <stdin>:2564:17, :2776:7
      Register_inst212 <= 32'h0;	// <stdin>:2564:17, :2777:7
      Register_inst213 <= 32'h0;	// <stdin>:2564:17, :2778:7
      Register_inst214 <= 32'h0;	// <stdin>:2564:17, :2779:7
      Register_inst215 <= 32'h0;	// <stdin>:2564:17, :2780:7
      Register_inst216 <= 32'h0;	// <stdin>:2564:17, :2781:7
      Register_inst217 <= 32'h0;	// <stdin>:2564:17, :2782:7
      Register_inst218 <= 32'h0;	// <stdin>:2564:17, :2783:7
      Register_inst219 <= 32'h0;	// <stdin>:2564:17, :2784:7
      Register_inst220 <= 32'h0;	// <stdin>:2564:17, :2785:7
      Register_inst221 <= 32'h0;	// <stdin>:2564:17, :2786:7
      Register_inst222 <= 32'h0;	// <stdin>:2564:17, :2787:7
      Register_inst223 <= 32'h0;	// <stdin>:2564:17, :2788:7
      Register_inst224 <= 32'h0;	// <stdin>:2564:17, :2789:7
      Register_inst225 <= 32'h0;	// <stdin>:2564:17, :2790:7
      Register_inst226 <= 32'h0;	// <stdin>:2564:17, :2791:7
      Register_inst227 <= 32'h0;	// <stdin>:2564:17, :2792:7
      Register_inst228 <= 32'h0;	// <stdin>:2564:17, :2793:7
      Register_inst229 <= 32'h0;	// <stdin>:2564:17, :2794:7
      Register_inst230 <= 32'h0;	// <stdin>:2564:17, :2795:7
      Register_inst231 <= 32'h0;	// <stdin>:2564:17, :2796:7
      Register_inst232 <= 32'h0;	// <stdin>:2564:17, :2797:7
      Register_inst233 <= 32'h0;	// <stdin>:2564:17, :2798:7
      Register_inst234 <= 32'h0;	// <stdin>:2564:17, :2799:7
      Register_inst235 <= 32'h0;	// <stdin>:2564:17, :2800:7
      Register_inst236 <= 32'h0;	// <stdin>:2564:17, :2801:7
      Register_inst237 <= 32'h0;	// <stdin>:2564:17, :2802:7
      Register_inst238 <= 32'h0;	// <stdin>:2564:17, :2803:7
      Register_inst239 <= 32'h0;	// <stdin>:2564:17, :2804:7
      Register_inst240 <= 32'h0;	// <stdin>:2564:17, :2805:7
      Register_inst241 <= 32'h0;	// <stdin>:2564:17, :2806:7
      Register_inst242 <= 32'h0;	// <stdin>:2564:17, :2807:7
      Register_inst243 <= 32'h0;	// <stdin>:2564:17, :2808:7
      Register_inst244 <= 32'h0;	// <stdin>:2564:17, :2809:7
      Register_inst245 <= 32'h0;	// <stdin>:2564:17, :2810:7
      Register_inst246 <= 32'h0;	// <stdin>:2564:17, :2811:7
      Register_inst247 <= 32'h0;	// <stdin>:2564:17, :2812:7
      Register_inst248 <= 32'h0;	// <stdin>:2564:17, :2813:7
      Register_inst249 <= 32'h0;	// <stdin>:2564:17, :2814:7
      Register_inst250 <= 32'h0;	// <stdin>:2564:17, :2815:7
      Register_inst251 <= 32'h0;	// <stdin>:2564:17, :2816:7
      Register_inst252 <= 32'h0;	// <stdin>:2564:17, :2817:7
      Register_inst253 <= 32'h0;	// <stdin>:2564:17, :2818:7
      Register_inst254 <= 32'h0;	// <stdin>:2564:17, :2819:7
      Register_inst255 <= 32'h0;	// <stdin>:2564:17, :2820:7
    end
    else begin	// <stdin>:2306:5
      Register_inst0 <= _T_255;	// <stdin>:2307:7
      Register_inst1 <= _T_256;	// <stdin>:2308:7
      Register_inst2 <= _T_257;	// <stdin>:2309:7
      Register_inst3 <= _T_258;	// <stdin>:2310:7
      Register_inst4 <= _T_259;	// <stdin>:2311:7
      Register_inst5 <= _T_260;	// <stdin>:2312:7
      Register_inst6 <= _T_261;	// <stdin>:2313:7
      Register_inst7 <= _T_262;	// <stdin>:2314:7
      Register_inst8 <= _T_263;	// <stdin>:2315:7
      Register_inst9 <= _T_264;	// <stdin>:2316:7
      Register_inst10 <= _T_265;	// <stdin>:2317:7
      Register_inst11 <= _T_266;	// <stdin>:2318:7
      Register_inst12 <= _T_267;	// <stdin>:2319:7
      Register_inst13 <= _T_268;	// <stdin>:2320:7
      Register_inst14 <= _T_269;	// <stdin>:2321:7
      Register_inst15 <= _T_270;	// <stdin>:2322:7
      Register_inst16 <= _T_271;	// <stdin>:2323:7
      Register_inst17 <= _T_272;	// <stdin>:2324:7
      Register_inst18 <= _T_273;	// <stdin>:2325:7
      Register_inst19 <= _T_274;	// <stdin>:2326:7
      Register_inst20 <= _T_275;	// <stdin>:2327:7
      Register_inst21 <= _T_276;	// <stdin>:2328:7
      Register_inst22 <= _T_277;	// <stdin>:2329:7
      Register_inst23 <= _T_278;	// <stdin>:2330:7
      Register_inst24 <= _T_279;	// <stdin>:2331:7
      Register_inst25 <= _T_280;	// <stdin>:2332:7
      Register_inst26 <= _T_281;	// <stdin>:2333:7
      Register_inst27 <= _T_282;	// <stdin>:2334:7
      Register_inst28 <= _T_283;	// <stdin>:2335:7
      Register_inst29 <= _T_284;	// <stdin>:2336:7
      Register_inst30 <= _T_285;	// <stdin>:2337:7
      Register_inst31 <= _T_286;	// <stdin>:2338:7
      Register_inst32 <= _T_287;	// <stdin>:2339:7
      Register_inst33 <= _T_288;	// <stdin>:2340:7
      Register_inst34 <= _T_289;	// <stdin>:2341:7
      Register_inst35 <= _T_290;	// <stdin>:2342:7
      Register_inst36 <= _T_291;	// <stdin>:2343:7
      Register_inst37 <= _T_292;	// <stdin>:2344:7
      Register_inst38 <= _T_293;	// <stdin>:2345:7
      Register_inst39 <= _T_294;	// <stdin>:2346:7
      Register_inst40 <= _T_295;	// <stdin>:2347:7
      Register_inst41 <= _T_296;	// <stdin>:2348:7
      Register_inst42 <= _T_297;	// <stdin>:2349:7
      Register_inst43 <= _T_298;	// <stdin>:2350:7
      Register_inst44 <= _T_299;	// <stdin>:2351:7
      Register_inst45 <= _T_300;	// <stdin>:2352:7
      Register_inst46 <= _T_301;	// <stdin>:2353:7
      Register_inst47 <= _T_302;	// <stdin>:2354:7
      Register_inst48 <= _T_303;	// <stdin>:2355:7
      Register_inst49 <= _T_304;	// <stdin>:2356:7
      Register_inst50 <= _T_305;	// <stdin>:2357:7
      Register_inst51 <= _T_306;	// <stdin>:2358:7
      Register_inst52 <= _T_307;	// <stdin>:2359:7
      Register_inst53 <= _T_308;	// <stdin>:2360:7
      Register_inst54 <= _T_309;	// <stdin>:2361:7
      Register_inst55 <= _T_310;	// <stdin>:2362:7
      Register_inst56 <= _T_311;	// <stdin>:2363:7
      Register_inst57 <= _T_312;	// <stdin>:2364:7
      Register_inst58 <= _T_313;	// <stdin>:2365:7
      Register_inst59 <= _T_314;	// <stdin>:2366:7
      Register_inst60 <= _T_315;	// <stdin>:2367:7
      Register_inst61 <= _T_316;	// <stdin>:2368:7
      Register_inst62 <= _T_317;	// <stdin>:2369:7
      Register_inst63 <= _T_318;	// <stdin>:2370:7
      Register_inst64 <= _T_319;	// <stdin>:2371:7
      Register_inst65 <= _T_320;	// <stdin>:2372:7
      Register_inst66 <= _T_321;	// <stdin>:2373:7
      Register_inst67 <= _T_322;	// <stdin>:2374:7
      Register_inst68 <= _T_323;	// <stdin>:2375:7
      Register_inst69 <= _T_324;	// <stdin>:2376:7
      Register_inst70 <= _T_325;	// <stdin>:2377:7
      Register_inst71 <= _T_326;	// <stdin>:2378:7
      Register_inst72 <= _T_327;	// <stdin>:2379:7
      Register_inst73 <= _T_328;	// <stdin>:2380:7
      Register_inst74 <= _T_329;	// <stdin>:2381:7
      Register_inst75 <= _T_330;	// <stdin>:2382:7
      Register_inst76 <= _T_331;	// <stdin>:2383:7
      Register_inst77 <= _T_332;	// <stdin>:2384:7
      Register_inst78 <= _T_333;	// <stdin>:2385:7
      Register_inst79 <= _T_334;	// <stdin>:2386:7
      Register_inst80 <= _T_335;	// <stdin>:2387:7
      Register_inst81 <= _T_336;	// <stdin>:2388:7
      Register_inst82 <= _T_337;	// <stdin>:2389:7
      Register_inst83 <= _T_338;	// <stdin>:2390:7
      Register_inst84 <= _T_339;	// <stdin>:2391:7
      Register_inst85 <= _T_340;	// <stdin>:2392:7
      Register_inst86 <= _T_341;	// <stdin>:2393:7
      Register_inst87 <= _T_342;	// <stdin>:2394:7
      Register_inst88 <= _T_343;	// <stdin>:2395:7
      Register_inst89 <= _T_344;	// <stdin>:2396:7
      Register_inst90 <= _T_345;	// <stdin>:2397:7
      Register_inst91 <= _T_346;	// <stdin>:2398:7
      Register_inst92 <= _T_347;	// <stdin>:2399:7
      Register_inst93 <= _T_348;	// <stdin>:2400:7
      Register_inst94 <= _T_349;	// <stdin>:2401:7
      Register_inst95 <= _T_350;	// <stdin>:2402:7
      Register_inst96 <= _T_351;	// <stdin>:2403:7
      Register_inst97 <= _T_352;	// <stdin>:2404:7
      Register_inst98 <= _T_353;	// <stdin>:2405:7
      Register_inst99 <= _T_354;	// <stdin>:2406:7
      Register_inst100 <= _T_355;	// <stdin>:2407:7
      Register_inst101 <= _T_356;	// <stdin>:2408:7
      Register_inst102 <= _T_357;	// <stdin>:2409:7
      Register_inst103 <= _T_358;	// <stdin>:2410:7
      Register_inst104 <= _T_359;	// <stdin>:2411:7
      Register_inst105 <= _T_360;	// <stdin>:2412:7
      Register_inst106 <= _T_361;	// <stdin>:2413:7
      Register_inst107 <= _T_362;	// <stdin>:2414:7
      Register_inst108 <= _T_363;	// <stdin>:2415:7
      Register_inst109 <= _T_364;	// <stdin>:2416:7
      Register_inst110 <= _T_365;	// <stdin>:2417:7
      Register_inst111 <= _T_366;	// <stdin>:2418:7
      Register_inst112 <= _T_367;	// <stdin>:2419:7
      Register_inst113 <= _T_368;	// <stdin>:2420:7
      Register_inst114 <= _T_369;	// <stdin>:2421:7
      Register_inst115 <= _T_370;	// <stdin>:2422:7
      Register_inst116 <= _T_371;	// <stdin>:2423:7
      Register_inst117 <= _T_372;	// <stdin>:2424:7
      Register_inst118 <= _T_373;	// <stdin>:2425:7
      Register_inst119 <= _T_374;	// <stdin>:2426:7
      Register_inst120 <= _T_375;	// <stdin>:2427:7
      Register_inst121 <= _T_376;	// <stdin>:2428:7
      Register_inst122 <= _T_377;	// <stdin>:2429:7
      Register_inst123 <= _T_378;	// <stdin>:2430:7
      Register_inst124 <= _T_379;	// <stdin>:2431:7
      Register_inst125 <= _T_380;	// <stdin>:2432:7
      Register_inst126 <= _T_381;	// <stdin>:2433:7
      Register_inst127 <= _T_382;	// <stdin>:2434:7
      Register_inst128 <= _T_383;	// <stdin>:2435:7
      Register_inst129 <= _T_384;	// <stdin>:2436:7
      Register_inst130 <= _T_385;	// <stdin>:2437:7
      Register_inst131 <= _T_386;	// <stdin>:2438:7
      Register_inst132 <= _T_387;	// <stdin>:2439:7
      Register_inst133 <= _T_388;	// <stdin>:2440:7
      Register_inst134 <= _T_389;	// <stdin>:2441:7
      Register_inst135 <= _T_390;	// <stdin>:2442:7
      Register_inst136 <= _T_391;	// <stdin>:2443:7
      Register_inst137 <= _T_392;	// <stdin>:2444:7
      Register_inst138 <= _T_393;	// <stdin>:2445:7
      Register_inst139 <= _T_394;	// <stdin>:2446:7
      Register_inst140 <= _T_395;	// <stdin>:2447:7
      Register_inst141 <= _T_396;	// <stdin>:2448:7
      Register_inst142 <= _T_397;	// <stdin>:2449:7
      Register_inst143 <= _T_398;	// <stdin>:2450:7
      Register_inst144 <= _T_399;	// <stdin>:2451:7
      Register_inst145 <= _T_400;	// <stdin>:2452:7
      Register_inst146 <= _T_401;	// <stdin>:2453:7
      Register_inst147 <= _T_402;	// <stdin>:2454:7
      Register_inst148 <= _T_403;	// <stdin>:2455:7
      Register_inst149 <= _T_404;	// <stdin>:2456:7
      Register_inst150 <= _T_405;	// <stdin>:2457:7
      Register_inst151 <= _T_406;	// <stdin>:2458:7
      Register_inst152 <= _T_407;	// <stdin>:2459:7
      Register_inst153 <= _T_408;	// <stdin>:2460:7
      Register_inst154 <= _T_409;	// <stdin>:2461:7
      Register_inst155 <= _T_410;	// <stdin>:2462:7
      Register_inst156 <= _T_411;	// <stdin>:2463:7
      Register_inst157 <= _T_412;	// <stdin>:2464:7
      Register_inst158 <= _T_413;	// <stdin>:2465:7
      Register_inst159 <= _T_414;	// <stdin>:2466:7
      Register_inst160 <= _T_415;	// <stdin>:2467:7
      Register_inst161 <= _T_416;	// <stdin>:2468:7
      Register_inst162 <= _T_417;	// <stdin>:2469:7
      Register_inst163 <= _T_418;	// <stdin>:2470:7
      Register_inst164 <= _T_419;	// <stdin>:2471:7
      Register_inst165 <= _T_420;	// <stdin>:2472:7
      Register_inst166 <= _T_421;	// <stdin>:2473:7
      Register_inst167 <= _T_422;	// <stdin>:2474:7
      Register_inst168 <= _T_423;	// <stdin>:2475:7
      Register_inst169 <= _T_424;	// <stdin>:2476:7
      Register_inst170 <= _T_425;	// <stdin>:2477:7
      Register_inst171 <= _T_426;	// <stdin>:2478:7
      Register_inst172 <= _T_427;	// <stdin>:2479:7
      Register_inst173 <= _T_428;	// <stdin>:2480:7
      Register_inst174 <= _T_429;	// <stdin>:2481:7
      Register_inst175 <= _T_430;	// <stdin>:2482:7
      Register_inst176 <= _T_431;	// <stdin>:2483:7
      Register_inst177 <= _T_432;	// <stdin>:2484:7
      Register_inst178 <= _T_433;	// <stdin>:2485:7
      Register_inst179 <= _T_434;	// <stdin>:2486:7
      Register_inst180 <= _T_435;	// <stdin>:2487:7
      Register_inst181 <= _T_436;	// <stdin>:2488:7
      Register_inst182 <= _T_437;	// <stdin>:2489:7
      Register_inst183 <= _T_438;	// <stdin>:2490:7
      Register_inst184 <= _T_439;	// <stdin>:2491:7
      Register_inst185 <= _T_440;	// <stdin>:2492:7
      Register_inst186 <= _T_441;	// <stdin>:2493:7
      Register_inst187 <= _T_442;	// <stdin>:2494:7
      Register_inst188 <= _T_443;	// <stdin>:2495:7
      Register_inst189 <= _T_444;	// <stdin>:2496:7
      Register_inst190 <= _T_445;	// <stdin>:2497:7
      Register_inst191 <= _T_446;	// <stdin>:2498:7
      Register_inst192 <= _T_447;	// <stdin>:2499:7
      Register_inst193 <= _T_448;	// <stdin>:2500:7
      Register_inst194 <= _T_449;	// <stdin>:2501:7
      Register_inst195 <= _T_450;	// <stdin>:2502:7
      Register_inst196 <= _T_451;	// <stdin>:2503:7
      Register_inst197 <= _T_452;	// <stdin>:2504:7
      Register_inst198 <= _T_453;	// <stdin>:2505:7
      Register_inst199 <= _T_454;	// <stdin>:2506:7
      Register_inst200 <= _T_455;	// <stdin>:2507:7
      Register_inst201 <= _T_456;	// <stdin>:2508:7
      Register_inst202 <= _T_457;	// <stdin>:2509:7
      Register_inst203 <= _T_458;	// <stdin>:2510:7
      Register_inst204 <= _T_459;	// <stdin>:2511:7
      Register_inst205 <= _T_460;	// <stdin>:2512:7
      Register_inst206 <= _T_461;	// <stdin>:2513:7
      Register_inst207 <= _T_462;	// <stdin>:2514:7
      Register_inst208 <= _T_463;	// <stdin>:2515:7
      Register_inst209 <= _T_464;	// <stdin>:2516:7
      Register_inst210 <= _T_465;	// <stdin>:2517:7
      Register_inst211 <= _T_466;	// <stdin>:2518:7
      Register_inst212 <= _T_467;	// <stdin>:2519:7
      Register_inst213 <= _T_468;	// <stdin>:2520:7
      Register_inst214 <= _T_469;	// <stdin>:2521:7
      Register_inst215 <= _T_470;	// <stdin>:2522:7
      Register_inst216 <= _T_471;	// <stdin>:2523:7
      Register_inst217 <= _T_472;	// <stdin>:2524:7
      Register_inst218 <= _T_473;	// <stdin>:2525:7
      Register_inst219 <= _T_474;	// <stdin>:2526:7
      Register_inst220 <= _T_475;	// <stdin>:2527:7
      Register_inst221 <= _T_476;	// <stdin>:2528:7
      Register_inst222 <= _T_477;	// <stdin>:2529:7
      Register_inst223 <= _T_478;	// <stdin>:2530:7
      Register_inst224 <= _T_479;	// <stdin>:2531:7
      Register_inst225 <= _T_480;	// <stdin>:2532:7
      Register_inst226 <= _T_481;	// <stdin>:2533:7
      Register_inst227 <= _T_482;	// <stdin>:2534:7
      Register_inst228 <= _T_483;	// <stdin>:2535:7
      Register_inst229 <= _T_484;	// <stdin>:2536:7
      Register_inst230 <= _T_485;	// <stdin>:2537:7
      Register_inst231 <= _T_486;	// <stdin>:2538:7
      Register_inst232 <= _T_487;	// <stdin>:2539:7
      Register_inst233 <= _T_488;	// <stdin>:2540:7
      Register_inst234 <= _T_489;	// <stdin>:2541:7
      Register_inst235 <= _T_490;	// <stdin>:2542:7
      Register_inst236 <= _T_491;	// <stdin>:2543:7
      Register_inst237 <= _T_492;	// <stdin>:2544:7
      Register_inst238 <= _T_493;	// <stdin>:2545:7
      Register_inst239 <= _T_494;	// <stdin>:2546:7
      Register_inst240 <= _T_495;	// <stdin>:2547:7
      Register_inst241 <= _T_496;	// <stdin>:2548:7
      Register_inst242 <= _T_497;	// <stdin>:2549:7
      Register_inst243 <= _T_498;	// <stdin>:2550:7
      Register_inst244 <= _T_499;	// <stdin>:2551:7
      Register_inst245 <= _T_500;	// <stdin>:2552:7
      Register_inst246 <= _T_501;	// <stdin>:2553:7
      Register_inst247 <= _T_502;	// <stdin>:2554:7
      Register_inst248 <= _T_503;	// <stdin>:2555:7
      Register_inst249 <= _T_504;	// <stdin>:2556:7
      Register_inst250 <= _T_505;	// <stdin>:2557:7
      Register_inst251 <= _T_506;	// <stdin>:2558:7
      Register_inst252 <= _T_507;	// <stdin>:2559:7
      Register_inst253 <= _T_508;	// <stdin>:2560:7
      Register_inst254 <= _T_509;	// <stdin>:2561:7
      Register_inst255 <= _T_510;	// <stdin>:2562:7
    end
  end // always @(posedge or posedge)
  initial begin	// <stdin>:2822:5
    Register_inst0 = 32'h0;	// <stdin>:2823:17, :2824:7
    Register_inst1 = 32'h0;	// <stdin>:2823:17, :2825:7
    Register_inst2 = 32'h0;	// <stdin>:2823:17, :2826:7
    Register_inst3 = 32'h0;	// <stdin>:2823:17, :2827:7
    Register_inst4 = 32'h0;	// <stdin>:2823:17, :2828:7
    Register_inst5 = 32'h0;	// <stdin>:2823:17, :2829:7
    Register_inst6 = 32'h0;	// <stdin>:2823:17, :2830:7
    Register_inst7 = 32'h0;	// <stdin>:2823:17, :2831:7
    Register_inst8 = 32'h0;	// <stdin>:2823:17, :2832:7
    Register_inst9 = 32'h0;	// <stdin>:2823:17, :2833:7
    Register_inst10 = 32'h0;	// <stdin>:2823:17, :2834:7
    Register_inst11 = 32'h0;	// <stdin>:2823:17, :2835:7
    Register_inst12 = 32'h0;	// <stdin>:2823:17, :2836:7
    Register_inst13 = 32'h0;	// <stdin>:2823:17, :2837:7
    Register_inst14 = 32'h0;	// <stdin>:2823:17, :2838:7
    Register_inst15 = 32'h0;	// <stdin>:2823:17, :2839:7
    Register_inst16 = 32'h0;	// <stdin>:2823:17, :2840:7
    Register_inst17 = 32'h0;	// <stdin>:2823:17, :2841:7
    Register_inst18 = 32'h0;	// <stdin>:2823:17, :2842:7
    Register_inst19 = 32'h0;	// <stdin>:2823:17, :2843:7
    Register_inst20 = 32'h0;	// <stdin>:2823:17, :2844:7
    Register_inst21 = 32'h0;	// <stdin>:2823:17, :2845:7
    Register_inst22 = 32'h0;	// <stdin>:2823:17, :2846:7
    Register_inst23 = 32'h0;	// <stdin>:2823:17, :2847:7
    Register_inst24 = 32'h0;	// <stdin>:2823:17, :2848:7
    Register_inst25 = 32'h0;	// <stdin>:2823:17, :2849:7
    Register_inst26 = 32'h0;	// <stdin>:2823:17, :2850:7
    Register_inst27 = 32'h0;	// <stdin>:2823:17, :2851:7
    Register_inst28 = 32'h0;	// <stdin>:2823:17, :2852:7
    Register_inst29 = 32'h0;	// <stdin>:2823:17, :2853:7
    Register_inst30 = 32'h0;	// <stdin>:2823:17, :2854:7
    Register_inst31 = 32'h0;	// <stdin>:2823:17, :2855:7
    Register_inst32 = 32'h0;	// <stdin>:2823:17, :2856:7
    Register_inst33 = 32'h0;	// <stdin>:2823:17, :2857:7
    Register_inst34 = 32'h0;	// <stdin>:2823:17, :2858:7
    Register_inst35 = 32'h0;	// <stdin>:2823:17, :2859:7
    Register_inst36 = 32'h0;	// <stdin>:2823:17, :2860:7
    Register_inst37 = 32'h0;	// <stdin>:2823:17, :2861:7
    Register_inst38 = 32'h0;	// <stdin>:2823:17, :2862:7
    Register_inst39 = 32'h0;	// <stdin>:2823:17, :2863:7
    Register_inst40 = 32'h0;	// <stdin>:2823:17, :2864:7
    Register_inst41 = 32'h0;	// <stdin>:2823:17, :2865:7
    Register_inst42 = 32'h0;	// <stdin>:2823:17, :2866:7
    Register_inst43 = 32'h0;	// <stdin>:2823:17, :2867:7
    Register_inst44 = 32'h0;	// <stdin>:2823:17, :2868:7
    Register_inst45 = 32'h0;	// <stdin>:2823:17, :2869:7
    Register_inst46 = 32'h0;	// <stdin>:2823:17, :2870:7
    Register_inst47 = 32'h0;	// <stdin>:2823:17, :2871:7
    Register_inst48 = 32'h0;	// <stdin>:2823:17, :2872:7
    Register_inst49 = 32'h0;	// <stdin>:2823:17, :2873:7
    Register_inst50 = 32'h0;	// <stdin>:2823:17, :2874:7
    Register_inst51 = 32'h0;	// <stdin>:2823:17, :2875:7
    Register_inst52 = 32'h0;	// <stdin>:2823:17, :2876:7
    Register_inst53 = 32'h0;	// <stdin>:2823:17, :2877:7
    Register_inst54 = 32'h0;	// <stdin>:2823:17, :2878:7
    Register_inst55 = 32'h0;	// <stdin>:2823:17, :2879:7
    Register_inst56 = 32'h0;	// <stdin>:2823:17, :2880:7
    Register_inst57 = 32'h0;	// <stdin>:2823:17, :2881:7
    Register_inst58 = 32'h0;	// <stdin>:2823:17, :2882:7
    Register_inst59 = 32'h0;	// <stdin>:2823:17, :2883:7
    Register_inst60 = 32'h0;	// <stdin>:2823:17, :2884:7
    Register_inst61 = 32'h0;	// <stdin>:2823:17, :2885:7
    Register_inst62 = 32'h0;	// <stdin>:2823:17, :2886:7
    Register_inst63 = 32'h0;	// <stdin>:2823:17, :2887:7
    Register_inst64 = 32'h0;	// <stdin>:2823:17, :2888:7
    Register_inst65 = 32'h0;	// <stdin>:2823:17, :2889:7
    Register_inst66 = 32'h0;	// <stdin>:2823:17, :2890:7
    Register_inst67 = 32'h0;	// <stdin>:2823:17, :2891:7
    Register_inst68 = 32'h0;	// <stdin>:2823:17, :2892:7
    Register_inst69 = 32'h0;	// <stdin>:2823:17, :2893:7
    Register_inst70 = 32'h0;	// <stdin>:2823:17, :2894:7
    Register_inst71 = 32'h0;	// <stdin>:2823:17, :2895:7
    Register_inst72 = 32'h0;	// <stdin>:2823:17, :2896:7
    Register_inst73 = 32'h0;	// <stdin>:2823:17, :2897:7
    Register_inst74 = 32'h0;	// <stdin>:2823:17, :2898:7
    Register_inst75 = 32'h0;	// <stdin>:2823:17, :2899:7
    Register_inst76 = 32'h0;	// <stdin>:2823:17, :2900:7
    Register_inst77 = 32'h0;	// <stdin>:2823:17, :2901:7
    Register_inst78 = 32'h0;	// <stdin>:2823:17, :2902:7
    Register_inst79 = 32'h0;	// <stdin>:2823:17, :2903:7
    Register_inst80 = 32'h0;	// <stdin>:2823:17, :2904:7
    Register_inst81 = 32'h0;	// <stdin>:2823:17, :2905:7
    Register_inst82 = 32'h0;	// <stdin>:2823:17, :2906:7
    Register_inst83 = 32'h0;	// <stdin>:2823:17, :2907:7
    Register_inst84 = 32'h0;	// <stdin>:2823:17, :2908:7
    Register_inst85 = 32'h0;	// <stdin>:2823:17, :2909:7
    Register_inst86 = 32'h0;	// <stdin>:2823:17, :2910:7
    Register_inst87 = 32'h0;	// <stdin>:2823:17, :2911:7
    Register_inst88 = 32'h0;	// <stdin>:2823:17, :2912:7
    Register_inst89 = 32'h0;	// <stdin>:2823:17, :2913:7
    Register_inst90 = 32'h0;	// <stdin>:2823:17, :2914:7
    Register_inst91 = 32'h0;	// <stdin>:2823:17, :2915:7
    Register_inst92 = 32'h0;	// <stdin>:2823:17, :2916:7
    Register_inst93 = 32'h0;	// <stdin>:2823:17, :2917:7
    Register_inst94 = 32'h0;	// <stdin>:2823:17, :2918:7
    Register_inst95 = 32'h0;	// <stdin>:2823:17, :2919:7
    Register_inst96 = 32'h0;	// <stdin>:2823:17, :2920:7
    Register_inst97 = 32'h0;	// <stdin>:2823:17, :2921:7
    Register_inst98 = 32'h0;	// <stdin>:2823:17, :2922:7
    Register_inst99 = 32'h0;	// <stdin>:2823:17, :2923:7
    Register_inst100 = 32'h0;	// <stdin>:2823:17, :2924:7
    Register_inst101 = 32'h0;	// <stdin>:2823:17, :2925:7
    Register_inst102 = 32'h0;	// <stdin>:2823:17, :2926:7
    Register_inst103 = 32'h0;	// <stdin>:2823:17, :2927:7
    Register_inst104 = 32'h0;	// <stdin>:2823:17, :2928:7
    Register_inst105 = 32'h0;	// <stdin>:2823:17, :2929:7
    Register_inst106 = 32'h0;	// <stdin>:2823:17, :2930:7
    Register_inst107 = 32'h0;	// <stdin>:2823:17, :2931:7
    Register_inst108 = 32'h0;	// <stdin>:2823:17, :2932:7
    Register_inst109 = 32'h0;	// <stdin>:2823:17, :2933:7
    Register_inst110 = 32'h0;	// <stdin>:2823:17, :2934:7
    Register_inst111 = 32'h0;	// <stdin>:2823:17, :2935:7
    Register_inst112 = 32'h0;	// <stdin>:2823:17, :2936:7
    Register_inst113 = 32'h0;	// <stdin>:2823:17, :2937:7
    Register_inst114 = 32'h0;	// <stdin>:2823:17, :2938:7
    Register_inst115 = 32'h0;	// <stdin>:2823:17, :2939:7
    Register_inst116 = 32'h0;	// <stdin>:2823:17, :2940:7
    Register_inst117 = 32'h0;	// <stdin>:2823:17, :2941:7
    Register_inst118 = 32'h0;	// <stdin>:2823:17, :2942:7
    Register_inst119 = 32'h0;	// <stdin>:2823:17, :2943:7
    Register_inst120 = 32'h0;	// <stdin>:2823:17, :2944:7
    Register_inst121 = 32'h0;	// <stdin>:2823:17, :2945:7
    Register_inst122 = 32'h0;	// <stdin>:2823:17, :2946:7
    Register_inst123 = 32'h0;	// <stdin>:2823:17, :2947:7
    Register_inst124 = 32'h0;	// <stdin>:2823:17, :2948:7
    Register_inst125 = 32'h0;	// <stdin>:2823:17, :2949:7
    Register_inst126 = 32'h0;	// <stdin>:2823:17, :2950:7
    Register_inst127 = 32'h0;	// <stdin>:2823:17, :2951:7
    Register_inst128 = 32'h0;	// <stdin>:2823:17, :2952:7
    Register_inst129 = 32'h0;	// <stdin>:2823:17, :2953:7
    Register_inst130 = 32'h0;	// <stdin>:2823:17, :2954:7
    Register_inst131 = 32'h0;	// <stdin>:2823:17, :2955:7
    Register_inst132 = 32'h0;	// <stdin>:2823:17, :2956:7
    Register_inst133 = 32'h0;	// <stdin>:2823:17, :2957:7
    Register_inst134 = 32'h0;	// <stdin>:2823:17, :2958:7
    Register_inst135 = 32'h0;	// <stdin>:2823:17, :2959:7
    Register_inst136 = 32'h0;	// <stdin>:2823:17, :2960:7
    Register_inst137 = 32'h0;	// <stdin>:2823:17, :2961:7
    Register_inst138 = 32'h0;	// <stdin>:2823:17, :2962:7
    Register_inst139 = 32'h0;	// <stdin>:2823:17, :2963:7
    Register_inst140 = 32'h0;	// <stdin>:2823:17, :2964:7
    Register_inst141 = 32'h0;	// <stdin>:2823:17, :2965:7
    Register_inst142 = 32'h0;	// <stdin>:2823:17, :2966:7
    Register_inst143 = 32'h0;	// <stdin>:2823:17, :2967:7
    Register_inst144 = 32'h0;	// <stdin>:2823:17, :2968:7
    Register_inst145 = 32'h0;	// <stdin>:2823:17, :2969:7
    Register_inst146 = 32'h0;	// <stdin>:2823:17, :2970:7
    Register_inst147 = 32'h0;	// <stdin>:2823:17, :2971:7
    Register_inst148 = 32'h0;	// <stdin>:2823:17, :2972:7
    Register_inst149 = 32'h0;	// <stdin>:2823:17, :2973:7
    Register_inst150 = 32'h0;	// <stdin>:2823:17, :2974:7
    Register_inst151 = 32'h0;	// <stdin>:2823:17, :2975:7
    Register_inst152 = 32'h0;	// <stdin>:2823:17, :2976:7
    Register_inst153 = 32'h0;	// <stdin>:2823:17, :2977:7
    Register_inst154 = 32'h0;	// <stdin>:2823:17, :2978:7
    Register_inst155 = 32'h0;	// <stdin>:2823:17, :2979:7
    Register_inst156 = 32'h0;	// <stdin>:2823:17, :2980:7
    Register_inst157 = 32'h0;	// <stdin>:2823:17, :2981:7
    Register_inst158 = 32'h0;	// <stdin>:2823:17, :2982:7
    Register_inst159 = 32'h0;	// <stdin>:2823:17, :2983:7
    Register_inst160 = 32'h0;	// <stdin>:2823:17, :2984:7
    Register_inst161 = 32'h0;	// <stdin>:2823:17, :2985:7
    Register_inst162 = 32'h0;	// <stdin>:2823:17, :2986:7
    Register_inst163 = 32'h0;	// <stdin>:2823:17, :2987:7
    Register_inst164 = 32'h0;	// <stdin>:2823:17, :2988:7
    Register_inst165 = 32'h0;	// <stdin>:2823:17, :2989:7
    Register_inst166 = 32'h0;	// <stdin>:2823:17, :2990:7
    Register_inst167 = 32'h0;	// <stdin>:2823:17, :2991:7
    Register_inst168 = 32'h0;	// <stdin>:2823:17, :2992:7
    Register_inst169 = 32'h0;	// <stdin>:2823:17, :2993:7
    Register_inst170 = 32'h0;	// <stdin>:2823:17, :2994:7
    Register_inst171 = 32'h0;	// <stdin>:2823:17, :2995:7
    Register_inst172 = 32'h0;	// <stdin>:2823:17, :2996:7
    Register_inst173 = 32'h0;	// <stdin>:2823:17, :2997:7
    Register_inst174 = 32'h0;	// <stdin>:2823:17, :2998:7
    Register_inst175 = 32'h0;	// <stdin>:2823:17, :2999:7
    Register_inst176 = 32'h0;	// <stdin>:2823:17, :3000:7
    Register_inst177 = 32'h0;	// <stdin>:2823:17, :3001:7
    Register_inst178 = 32'h0;	// <stdin>:2823:17, :3002:7
    Register_inst179 = 32'h0;	// <stdin>:2823:17, :3003:7
    Register_inst180 = 32'h0;	// <stdin>:2823:17, :3004:7
    Register_inst181 = 32'h0;	// <stdin>:2823:17, :3005:7
    Register_inst182 = 32'h0;	// <stdin>:2823:17, :3006:7
    Register_inst183 = 32'h0;	// <stdin>:2823:17, :3007:7
    Register_inst184 = 32'h0;	// <stdin>:2823:17, :3008:7
    Register_inst185 = 32'h0;	// <stdin>:2823:17, :3009:7
    Register_inst186 = 32'h0;	// <stdin>:2823:17, :3010:7
    Register_inst187 = 32'h0;	// <stdin>:2823:17, :3011:7
    Register_inst188 = 32'h0;	// <stdin>:2823:17, :3012:7
    Register_inst189 = 32'h0;	// <stdin>:2823:17, :3013:7
    Register_inst190 = 32'h0;	// <stdin>:2823:17, :3014:7
    Register_inst191 = 32'h0;	// <stdin>:2823:17, :3015:7
    Register_inst192 = 32'h0;	// <stdin>:2823:17, :3016:7
    Register_inst193 = 32'h0;	// <stdin>:2823:17, :3017:7
    Register_inst194 = 32'h0;	// <stdin>:2823:17, :3018:7
    Register_inst195 = 32'h0;	// <stdin>:2823:17, :3019:7
    Register_inst196 = 32'h0;	// <stdin>:2823:17, :3020:7
    Register_inst197 = 32'h0;	// <stdin>:2823:17, :3021:7
    Register_inst198 = 32'h0;	// <stdin>:2823:17, :3022:7
    Register_inst199 = 32'h0;	// <stdin>:2823:17, :3023:7
    Register_inst200 = 32'h0;	// <stdin>:2823:17, :3024:7
    Register_inst201 = 32'h0;	// <stdin>:2823:17, :3025:7
    Register_inst202 = 32'h0;	// <stdin>:2823:17, :3026:7
    Register_inst203 = 32'h0;	// <stdin>:2823:17, :3027:7
    Register_inst204 = 32'h0;	// <stdin>:2823:17, :3028:7
    Register_inst205 = 32'h0;	// <stdin>:2823:17, :3029:7
    Register_inst206 = 32'h0;	// <stdin>:2823:17, :3030:7
    Register_inst207 = 32'h0;	// <stdin>:2823:17, :3031:7
    Register_inst208 = 32'h0;	// <stdin>:2823:17, :3032:7
    Register_inst209 = 32'h0;	// <stdin>:2823:17, :3033:7
    Register_inst210 = 32'h0;	// <stdin>:2823:17, :3034:7
    Register_inst211 = 32'h0;	// <stdin>:2823:17, :3035:7
    Register_inst212 = 32'h0;	// <stdin>:2823:17, :3036:7
    Register_inst213 = 32'h0;	// <stdin>:2823:17, :3037:7
    Register_inst214 = 32'h0;	// <stdin>:2823:17, :3038:7
    Register_inst215 = 32'h0;	// <stdin>:2823:17, :3039:7
    Register_inst216 = 32'h0;	// <stdin>:2823:17, :3040:7
    Register_inst217 = 32'h0;	// <stdin>:2823:17, :3041:7
    Register_inst218 = 32'h0;	// <stdin>:2823:17, :3042:7
    Register_inst219 = 32'h0;	// <stdin>:2823:17, :3043:7
    Register_inst220 = 32'h0;	// <stdin>:2823:17, :3044:7
    Register_inst221 = 32'h0;	// <stdin>:2823:17, :3045:7
    Register_inst222 = 32'h0;	// <stdin>:2823:17, :3046:7
    Register_inst223 = 32'h0;	// <stdin>:2823:17, :3047:7
    Register_inst224 = 32'h0;	// <stdin>:2823:17, :3048:7
    Register_inst225 = 32'h0;	// <stdin>:2823:17, :3049:7
    Register_inst226 = 32'h0;	// <stdin>:2823:17, :3050:7
    Register_inst227 = 32'h0;	// <stdin>:2823:17, :3051:7
    Register_inst228 = 32'h0;	// <stdin>:2823:17, :3052:7
    Register_inst229 = 32'h0;	// <stdin>:2823:17, :3053:7
    Register_inst230 = 32'h0;	// <stdin>:2823:17, :3054:7
    Register_inst231 = 32'h0;	// <stdin>:2823:17, :3055:7
    Register_inst232 = 32'h0;	// <stdin>:2823:17, :3056:7
    Register_inst233 = 32'h0;	// <stdin>:2823:17, :3057:7
    Register_inst234 = 32'h0;	// <stdin>:2823:17, :3058:7
    Register_inst235 = 32'h0;	// <stdin>:2823:17, :3059:7
    Register_inst236 = 32'h0;	// <stdin>:2823:17, :3060:7
    Register_inst237 = 32'h0;	// <stdin>:2823:17, :3061:7
    Register_inst238 = 32'h0;	// <stdin>:2823:17, :3062:7
    Register_inst239 = 32'h0;	// <stdin>:2823:17, :3063:7
    Register_inst240 = 32'h0;	// <stdin>:2823:17, :3064:7
    Register_inst241 = 32'h0;	// <stdin>:2823:17, :3065:7
    Register_inst242 = 32'h0;	// <stdin>:2823:17, :3066:7
    Register_inst243 = 32'h0;	// <stdin>:2823:17, :3067:7
    Register_inst244 = 32'h0;	// <stdin>:2823:17, :3068:7
    Register_inst245 = 32'h0;	// <stdin>:2823:17, :3069:7
    Register_inst246 = 32'h0;	// <stdin>:2823:17, :3070:7
    Register_inst247 = 32'h0;	// <stdin>:2823:17, :3071:7
    Register_inst248 = 32'h0;	// <stdin>:2823:17, :3072:7
    Register_inst249 = 32'h0;	// <stdin>:2823:17, :3073:7
    Register_inst250 = 32'h0;	// <stdin>:2823:17, :3074:7
    Register_inst251 = 32'h0;	// <stdin>:2823:17, :3075:7
    Register_inst252 = 32'h0;	// <stdin>:2823:17, :3076:7
    Register_inst253 = 32'h0;	// <stdin>:2823:17, :3077:7
    Register_inst254 = 32'h0;	// <stdin>:2823:17, :3078:7
    Register_inst255 = 32'h0;	// <stdin>:2823:17, :3079:7
  end // initial
  assign _T = Register_inst255;	// <stdin>:3081:13
  wire [255:0][31:0] _tmp_511 = {{_T_254}, {_T_253}, {_T_252}, {_T_251}, {_T_250}, {_T_249}, {_T_248}, {_T_247}, {_T_246}, {_T_245}, {_T_244}, {_T_243}, {_T_242}, {_T_241}, {_T_240}, {_T_239}, {_T_238}, {_T_237}, {_T_236}, {_T_235}, {_T_234}, {_T_233}, {_T_232}, {_T_231}, {_T_230}, {_T_229}, {_T_228}, {_T_227}, {_T_226}, {_T_225}, {_T_224}, {_T_223}, {_T_222}, {_T_221}, {_T_220}, {_T_219}, {_T_218}, {_T_217}, {_T_216}, {_T_215}, {_T_214}, {_T_213}, {_T_212}, {_T_211}, {_T_210}, {_T_209}, {_T_208}, {_T_207}, {_T_206}, {_T_205}, {_T_204}, {_T_203}, {_T_202}, {_T_201}, {_T_200}, {_T_199}, {_T_198}, {_T_197}, {_T_196}, {_T_195}, {_T_194}, {_T_193}, {_T_192}, {_T_191}, {_T_190}, {_T_189}, {_T_188}, {_T_187}, {_T_186}, {_T_185}, {_T_184}, {_T_183}, {_T_182}, {_T_181}, {_T_180}, {_T_179}, {_T_178}, {_T_177}, {_T_176}, {_T_175}, {_T_174}, {_T_173}, {_T_172}, {_T_171}, {_T_170}, {_T_169}, {_T_168}, {_T_167}, {_T_166}, {_T_165}, {_T_164}, {_T_163}, {_T_162}, {_T_161}, {_T_160}, {_T_159}, {_T_158}, {_T_157}, {_T_156}, {_T_155}, {_T_154}, {_T_153}, {_T_152}, {_T_151}, {_T_150}, {_T_149}, {_T_148}, {_T_147}, {_T_146}, {_T_145}, {_T_144}, {_T_143}, {_T_142}, {_T_141}, {_T_140}, {_T_139}, {_T_138}, {_T_137}, {_T_136}, {_T_135}, {_T_134}, {_T_133}, {_T_132}, {_T_131}, {_T_130}, {_T_129}, {_T_128}, {_T_127}, {_T_126}, {_T_125}, {_T_124}, {_T_123}, {_T_122}, {_T_121}, {_T_120}, {_T_119}, {_T_118}, {_T_117}, {_T_116}, {_T_115}, {_T_114}, {_T_113}, {_T_112}, {_T_111}, {_T_110}, {_T_109}, {_T_108}, {_T_107}, {_T_106}, {_T_105}, {_T_104}, {_T_103}, {_T_102}, {_T_101}, {_T_100}, {_T_99}, {_T_98}, {_T_97}, {_T_96}, {_T_95}, {_T_94}, {_T_93}, {_T_92}, {_T_91}, {_T_90}, {_T_89}, {_T_88}, {_T_87}, {_T_86}, {_T_85}, {_T_84}, {_T_83}, {_T_82}, {_T_81}, {_T_80}, {_T_79}, {_T_78}, {_T_77}, {_T_76}, {_T_75}, {_T_74}, {_T_73}, {_T_72}, {_T_71}, {_T_70}, {_T_69}, {_T_68}, {_T_67}, {_T_66}, {_T_65}, {_T_64}, {_T_63}, {_T_62}, {_T_61}, {_T_60}, {_T_59}, {_T_58}, {_T_57}, {_T_56}, {_T_55}, {_T_54}, {_T_53}, {_T_52}, {_T_51}, {_T_50}, {_T_49}, {_T_48}, {_T_47}, {_T_46}, {_T_45}, {_T_44}, {_T_43}, {_T_42}, {_T_41}, {_T_40}, {_T_39}, {_T_38}, {_T_37}, {_T_36}, {_T_35}, {_T_34}, {_T_33}, {_T_32}, {_T_31}, {_T_30}, {_T_29}, {_T_28}, {_T_27}, {_T_26}, {_T_25}, {_T_24}, {_T_23}, {_T_22}, {_T_21}, {_T_20}, {_T_19}, {_T_18}, {_T_17}, {_T_16}, {_T_15}, {_T_14}, {_T_13}, {_T_12}, {_T_11}, {_T_10}, {_T_9}, {_T_8}, {_T_7}, {_T_6}, {_T_5}, {_T_4}, {_T_3}, {_T_2}, {_T_1}, {_T_0}, {_T}};	// <stdin>:266:10, :274:11, :282:11, :290:11, :298:11, :306:11, :314:11, :322:11, :330:11, :338:11, :346:11, :354:11, :362:11, :370:11, :378:12, :386:12, :394:12, :402:12, :410:12, :418:12, :426:12, :434:12, :442:12, :450:12, :458:12, :466:12, :474:12, :482:12, :490:12, :498:12, :506:12, :514:12, :522:12, :530:12, :538:12, :546:12, :554:12, :562:12, :570:12, :578:12, :586:12, :594:12, :602:12, :610:12, :618:12, :626:12, :634:12, :642:12, :650:12, :658:12, :666:12, :674:12, :682:12, :690:12, :698:12, :706:12, :714:12, :722:12, :730:12, :738:12, :746:12, :754:12, :762:12, :770:12, :778:12, :786:12, :794:12, :802:12, :810:12, :818:12, :826:12, :834:12, :842:12, :850:12, :858:12, :866:12, :874:12, :882:12, :890:12, :898:12, :906:12, :914:12, :922:12, :930:12, :938:12, :946:12, :954:12, :962:12, :970:12, :978:12, :986:12, :994:12, :1002:12, :1010:12, :1018:12, :1026:12, :1034:12, :1042:12, :1050:12, :1058:12, :1066:12, :1074:12, :1082:12, :1090:12, :1098:12, :1106:12, :1114:12, :1122:12, :1130:12, :1138:12, :1146:12, :1154:12, :1162:12, :1170:12, :1178:12, :1186:12, :1194:12, :1202:12, :1210:12, :1218:12, :1226:12, :1234:12, :1242:12, :1250:12, :1258:12, :1266:12, :1274:12, :1282:12, :1290:12, :1298:12, :1306:12, :1314:12, :1322:12, :1330:12, :1338:12, :1346:12, :1354:12, :1362:12, :1370:12, :1378:12, :1386:12, :1394:12, :1402:13, :1410:13, :1418:13, :1426:13, :1434:13, :1442:13, :1450:13, :1458:13, :1466:13, :1474:13, :1482:13, :1490:13, :1498:13, :1506:13, :1514:13, :1522:13, :1530:13, :1538:13, :1546:13, :1554:13, :1562:13, :1570:13, :1578:13, :1586:13, :1594:13, :1602:13, :1610:13, :1618:13, :1626:13, :1634:13, :1642:13, :1650:13, :1658:13, :1666:13, :1674:13, :1682:13, :1690:13, :1698:13, :1706:13, :1714:13, :1722:13, :1730:13, :1738:13, :1746:13, :1754:13, :1762:13, :1770:13, :1778:13, :1786:13, :1794:13, :1802:13, :1810:13, :1818:13, :1826:13, :1834:13, :1842:13, :1850:13, :1858:13, :1866:13, :1874:13, :1882:13, :1890:13, :1898:13, :1906:13, :1914:13, :1922:13, :1930:13, :1938:13, :1946:13, :1954:13, :1962:13, :1970:13, :1978:13, :1986:13, :1994:13, :2002:13, :2010:13, :2018:13, :2026:13, :2034:13, :2042:13, :2050:13, :2058:13, :2066:13, :2074:13, :2082:13, :2090:13, :2098:13, :2106:13, :2114:13, :2122:13, :2130:13, :2138:13, :2146:13, :2154:13, :2162:13, :2170:13, :2178:13, :2186:13, :2194:13, :2202:13, :2210:13, :2218:13, :2226:13, :2234:13, :2242:13, :2250:13, :2258:13, :2266:13, :2274:13, :2282:13, :2290:13, :2298:13, :3081:13, :3084:13
  wire [255:0][31:0] _tmp = {{_T_254}, {_T_253}, {_T_252}, {_T_251}, {_T_250}, {_T_249}, {_T_248}, {_T_247}, {_T_246}, {_T_245}, {_T_244}, {_T_243}, {_T_242}, {_T_241}, {_T_240}, {_T_239}, {_T_238}, {_T_237}, {_T_236}, {_T_235}, {_T_234}, {_T_233}, {_T_232}, {_T_231}, {_T_230}, {_T_229}, {_T_228}, {_T_227}, {_T_226}, {_T_225}, {_T_224}, {_T_223}, {_T_222}, {_T_221}, {_T_220}, {_T_219}, {_T_218}, {_T_217}, {_T_216}, {_T_215}, {_T_214}, {_T_213}, {_T_212}, {_T_211}, {_T_210}, {_T_209}, {_T_208}, {_T_207}, {_T_206}, {_T_205}, {_T_204}, {_T_203}, {_T_202}, {_T_201}, {_T_200}, {_T_199}, {_T_198}, {_T_197}, {_T_196}, {_T_195}, {_T_194}, {_T_193}, {_T_192}, {_T_191}, {_T_190}, {_T_189}, {_T_188}, {_T_187}, {_T_186}, {_T_185}, {_T_184}, {_T_183}, {_T_182}, {_T_181}, {_T_180}, {_T_179}, {_T_178}, {_T_177}, {_T_176}, {_T_175}, {_T_174}, {_T_173}, {_T_172}, {_T_171}, {_T_170}, {_T_169}, {_T_168}, {_T_167}, {_T_166}, {_T_165}, {_T_164}, {_T_163}, {_T_162}, {_T_161}, {_T_160}, {_T_159}, {_T_158}, {_T_157}, {_T_156}, {_T_155}, {_T_154}, {_T_153}, {_T_152}, {_T_151}, {_T_150}, {_T_149}, {_T_148}, {_T_147}, {_T_146}, {_T_145}, {_T_144}, {_T_143}, {_T_142}, {_T_141}, {_T_140}, {_T_139}, {_T_138}, {_T_137}, {_T_136}, {_T_135}, {_T_134}, {_T_133}, {_T_132}, {_T_131}, {_T_130}, {_T_129}, {_T_128}, {_T_127}, {_T_126}, {_T_125}, {_T_124}, {_T_123}, {_T_122}, {_T_121}, {_T_120}, {_T_119}, {_T_118}, {_T_117}, {_T_116}, {_T_115}, {_T_114}, {_T_113}, {_T_112}, {_T_111}, {_T_110}, {_T_109}, {_T_108}, {_T_107}, {_T_106}, {_T_105}, {_T_104}, {_T_103}, {_T_102}, {_T_101}, {_T_100}, {_T_99}, {_T_98}, {_T_97}, {_T_96}, {_T_95}, {_T_94}, {_T_93}, {_T_92}, {_T_91}, {_T_90}, {_T_89}, {_T_88}, {_T_87}, {_T_86}, {_T_85}, {_T_84}, {_T_83}, {_T_82}, {_T_81}, {_T_80}, {_T_79}, {_T_78}, {_T_77}, {_T_76}, {_T_75}, {_T_74}, {_T_73}, {_T_72}, {_T_71}, {_T_70}, {_T_69}, {_T_68}, {_T_67}, {_T_66}, {_T_65}, {_T_64}, {_T_63}, {_T_62}, {_T_61}, {_T_60}, {_T_59}, {_T_58}, {_T_57}, {_T_56}, {_T_55}, {_T_54}, {_T_53}, {_T_52}, {_T_51}, {_T_50}, {_T_49}, {_T_48}, {_T_47}, {_T_46}, {_T_45}, {_T_44}, {_T_43}, {_T_42}, {_T_41}, {_T_40}, {_T_39}, {_T_38}, {_T_37}, {_T_36}, {_T_35}, {_T_34}, {_T_33}, {_T_32}, {_T_31}, {_T_30}, {_T_29}, {_T_28}, {_T_27}, {_T_26}, {_T_25}, {_T_24}, {_T_23}, {_T_22}, {_T_21}, {_T_20}, {_T_19}, {_T_18}, {_T_17}, {_T_16}, {_T_15}, {_T_14}, {_T_13}, {_T_12}, {_T_11}, {_T_10}, {_T_9}, {_T_8}, {_T_7}, {_T_6}, {_T_5}, {_T_4}, {_T_3}, {_T_2}, {_T_1}, {_T_0}, {_T}};	// <stdin>:266:10, :274:11, :282:11, :290:11, :298:11, :306:11, :314:11, :322:11, :330:11, :338:11, :346:11, :354:11, :362:11, :370:11, :378:12, :386:12, :394:12, :402:12, :410:12, :418:12, :426:12, :434:12, :442:12, :450:12, :458:12, :466:12, :474:12, :482:12, :490:12, :498:12, :506:12, :514:12, :522:12, :530:12, :538:12, :546:12, :554:12, :562:12, :570:12, :578:12, :586:12, :594:12, :602:12, :610:12, :618:12, :626:12, :634:12, :642:12, :650:12, :658:12, :666:12, :674:12, :682:12, :690:12, :698:12, :706:12, :714:12, :722:12, :730:12, :738:12, :746:12, :754:12, :762:12, :770:12, :778:12, :786:12, :794:12, :802:12, :810:12, :818:12, :826:12, :834:12, :842:12, :850:12, :858:12, :866:12, :874:12, :882:12, :890:12, :898:12, :906:12, :914:12, :922:12, :930:12, :938:12, :946:12, :954:12, :962:12, :970:12, :978:12, :986:12, :994:12, :1002:12, :1010:12, :1018:12, :1026:12, :1034:12, :1042:12, :1050:12, :1058:12, :1066:12, :1074:12, :1082:12, :1090:12, :1098:12, :1106:12, :1114:12, :1122:12, :1130:12, :1138:12, :1146:12, :1154:12, :1162:12, :1170:12, :1178:12, :1186:12, :1194:12, :1202:12, :1210:12, :1218:12, :1226:12, :1234:12, :1242:12, :1250:12, :1258:12, :1266:12, :1274:12, :1282:12, :1290:12, :1298:12, :1306:12, :1314:12, :1322:12, :1330:12, :1338:12, :1346:12, :1354:12, :1362:12, :1370:12, :1378:12, :1386:12, :1394:12, :1402:13, :1410:13, :1418:13, :1426:13, :1434:13, :1442:13, :1450:13, :1458:13, :1466:13, :1474:13, :1482:13, :1490:13, :1498:13, :1506:13, :1514:13, :1522:13, :1530:13, :1538:13, :1546:13, :1554:13, :1562:13, :1570:13, :1578:13, :1586:13, :1594:13, :1602:13, :1610:13, :1618:13, :1626:13, :1634:13, :1642:13, :1650:13, :1658:13, :1666:13, :1674:13, :1682:13, :1690:13, :1698:13, :1706:13, :1714:13, :1722:13, :1730:13, :1738:13, :1746:13, :1754:13, :1762:13, :1770:13, :1778:13, :1786:13, :1794:13, :1802:13, :1810:13, :1818:13, :1826:13, :1834:13, :1842:13, :1850:13, :1858:13, :1866:13, :1874:13, :1882:13, :1890:13, :1898:13, :1906:13, :1914:13, :1922:13, :1930:13, :1938:13, :1946:13, :1954:13, :1962:13, :1970:13, :1978:13, :1986:13, :1994:13, :2002:13, :2010:13, :2018:13, :2026:13, :2034:13, :2042:13, :2050:13, :2058:13, :2066:13, :2074:13, :2082:13, :2090:13, :2098:13, :2106:13, :2114:13, :2122:13, :2130:13, :2138:13, :2146:13, :2154:13, :2162:13, :2170:13, :2178:13, :2186:13, :2194:13, :2202:13, :2210:13, :2218:13, :2226:13, :2234:13, :2242:13, :2250:13, :2258:13, :2266:13, :2274:13, :2282:13, :2290:13, :2298:13, :3081:13, :3082:13
  assign file_read_0_data = _tmp[file_read_0_addr];	// <stdin>:266:10, :274:11, :282:11, :290:11, :298:11, :306:11, :314:11, :322:11, :330:11, :338:11, :346:11, :354:11, :362:11, :370:11, :378:12, :386:12, :394:12, :402:12, :410:12, :418:12, :426:12, :434:12, :442:12, :450:12, :458:12, :466:12, :474:12, :482:12, :490:12, :498:12, :506:12, :514:12, :522:12, :530:12, :538:12, :546:12, :554:12, :562:12, :570:12, :578:12, :586:12, :594:12, :602:12, :610:12, :618:12, :626:12, :634:12, :642:12, :650:12, :658:12, :666:12, :674:12, :682:12, :690:12, :698:12, :706:12, :714:12, :722:12, :730:12, :738:12, :746:12, :754:12, :762:12, :770:12, :778:12, :786:12, :794:12, :802:12, :810:12, :818:12, :826:12, :834:12, :842:12, :850:12, :858:12, :866:12, :874:12, :882:12, :890:12, :898:12, :906:12, :914:12, :922:12, :930:12, :938:12, :946:12, :954:12, :962:12, :970:12, :978:12, :986:12, :994:12, :1002:12, :1010:12, :1018:12, :1026:12, :1034:12, :1042:12, :1050:12, :1058:12, :1066:12, :1074:12, :1082:12, :1090:12, :1098:12, :1106:12, :1114:12, :1122:12, :1130:12, :1138:12, :1146:12, :1154:12, :1162:12, :1170:12, :1178:12, :1186:12, :1194:12, :1202:12, :1210:12, :1218:12, :1226:12, :1234:12, :1242:12, :1250:12, :1258:12, :1266:12, :1274:12, :1282:12, :1290:12, :1298:12, :1306:12, :1314:12, :1322:12, :1330:12, :1338:12, :1346:12, :1354:12, :1362:12, :1370:12, :1378:12, :1386:12, :1394:12, :1402:13, :1410:13, :1418:13, :1426:13, :1434:13, :1442:13, :1450:13, :1458:13, :1466:13, :1474:13, :1482:13, :1490:13, :1498:13, :1506:13, :1514:13, :1522:13, :1530:13, :1538:13, :1546:13, :1554:13, :1562:13, :1570:13, :1578:13, :1586:13, :1594:13, :1602:13, :1610:13, :1618:13, :1626:13, :1634:13, :1642:13, :1650:13, :1658:13, :1666:13, :1674:13, :1682:13, :1690:13, :1698:13, :1706:13, :1714:13, :1722:13, :1730:13, :1738:13, :1746:13, :1754:13, :1762:13, :1770:13, :1778:13, :1786:13, :1794:13, :1802:13, :1810:13, :1818:13, :1826:13, :1834:13, :1842:13, :1850:13, :1858:13, :1866:13, :1874:13, :1882:13, :1890:13, :1898:13, :1906:13, :1914:13, :1922:13, :1930:13, :1938:13, :1946:13, :1954:13, :1962:13, :1970:13, :1978:13, :1986:13, :1994:13, :2002:13, :2010:13, :2018:13, :2026:13, :2034:13, :2042:13, :2050:13, :2058:13, :2066:13, :2074:13, :2082:13, :2090:13, :2098:13, :2106:13, :2114:13, :2122:13, :2130:13, :2138:13, :2146:13, :2154:13, :2162:13, :2170:13, :2178:13, :2186:13, :2194:13, :2202:13, :2210:13, :2218:13, :2226:13, :2234:13, :2242:13, :2250:13, :2258:13, :2266:13, :2274:13, :2282:13, :2290:13, :2298:13, :3081:13, :3083:13, :3086:5
  assign file_read_1_data = _tmp_511[file_read_1_addr];	// <stdin>:266:10, :274:11, :282:11, :290:11, :298:11, :306:11, :314:11, :322:11, :330:11, :338:11, :346:11, :354:11, :362:11, :370:11, :378:12, :386:12, :394:12, :402:12, :410:12, :418:12, :426:12, :434:12, :442:12, :450:12, :458:12, :466:12, :474:12, :482:12, :490:12, :498:12, :506:12, :514:12, :522:12, :530:12, :538:12, :546:12, :554:12, :562:12, :570:12, :578:12, :586:12, :594:12, :602:12, :610:12, :618:12, :626:12, :634:12, :642:12, :650:12, :658:12, :666:12, :674:12, :682:12, :690:12, :698:12, :706:12, :714:12, :722:12, :730:12, :738:12, :746:12, :754:12, :762:12, :770:12, :778:12, :786:12, :794:12, :802:12, :810:12, :818:12, :826:12, :834:12, :842:12, :850:12, :858:12, :866:12, :874:12, :882:12, :890:12, :898:12, :906:12, :914:12, :922:12, :930:12, :938:12, :946:12, :954:12, :962:12, :970:12, :978:12, :986:12, :994:12, :1002:12, :1010:12, :1018:12, :1026:12, :1034:12, :1042:12, :1050:12, :1058:12, :1066:12, :1074:12, :1082:12, :1090:12, :1098:12, :1106:12, :1114:12, :1122:12, :1130:12, :1138:12, :1146:12, :1154:12, :1162:12, :1170:12, :1178:12, :1186:12, :1194:12, :1202:12, :1210:12, :1218:12, :1226:12, :1234:12, :1242:12, :1250:12, :1258:12, :1266:12, :1274:12, :1282:12, :1290:12, :1298:12, :1306:12, :1314:12, :1322:12, :1330:12, :1338:12, :1346:12, :1354:12, :1362:12, :1370:12, :1378:12, :1386:12, :1394:12, :1402:13, :1410:13, :1418:13, :1426:13, :1434:13, :1442:13, :1450:13, :1458:13, :1466:13, :1474:13, :1482:13, :1490:13, :1498:13, :1506:13, :1514:13, :1522:13, :1530:13, :1538:13, :1546:13, :1554:13, :1562:13, :1570:13, :1578:13, :1586:13, :1594:13, :1602:13, :1610:13, :1618:13, :1626:13, :1634:13, :1642:13, :1650:13, :1658:13, :1666:13, :1674:13, :1682:13, :1690:13, :1698:13, :1706:13, :1714:13, :1722:13, :1730:13, :1738:13, :1746:13, :1754:13, :1762:13, :1770:13, :1778:13, :1786:13, :1794:13, :1802:13, :1810:13, :1818:13, :1826:13, :1834:13, :1842:13, :1850:13, :1858:13, :1866:13, :1874:13, :1882:13, :1890:13, :1898:13, :1906:13, :1914:13, :1922:13, :1930:13, :1938:13, :1946:13, :1954:13, :1962:13, :1970:13, :1978:13, :1986:13, :1994:13, :2002:13, :2010:13, :2018:13, :2026:13, :2034:13, :2042:13, :2050:13, :2058:13, :2066:13, :2074:13, :2082:13, :2090:13, :2098:13, :2106:13, :2114:13, :2122:13, :2130:13, :2138:13, :2146:13, :2154:13, :2162:13, :2170:13, :2178:13, :2186:13, :2194:13, :2202:13, :2210:13, :2218:13, :2226:13, :2234:13, :2242:13, :2250:13, :2258:13, :2266:13, :2274:13, :2282:13, :2290:13, :2298:13, :3081:13, :3085:13, :3086:5
endmodule

module code(
  input                                                        CLK, ASYNCRESET,
  input  [7:0]                                                 code_read_0_addr,
  input  struct packed {logic [31:0] data; logic [7:0] addr; } write_0,
  input                                                        write_0_en,
  output [31:0]                                                code_read_0_data);

  wire [31:0] _T;	// <stdin>:6167:13
  wire [31:0] _T_0;	// <stdin>:5384:13
  wire [31:0] _T_1;	// <stdin>:5376:13
  wire [31:0] _T_2;	// <stdin>:5368:13
  wire [31:0] _T_3;	// <stdin>:5360:13
  wire [31:0] _T_4;	// <stdin>:5352:13
  wire [31:0] _T_5;	// <stdin>:5344:13
  wire [31:0] _T_6;	// <stdin>:5336:13
  wire [31:0] _T_7;	// <stdin>:5328:13
  wire [31:0] _T_8;	// <stdin>:5320:13
  wire [31:0] _T_9;	// <stdin>:5312:13
  wire [31:0] _T_10;	// <stdin>:5304:13
  wire [31:0] _T_11;	// <stdin>:5296:13
  wire [31:0] _T_12;	// <stdin>:5288:13
  wire [31:0] _T_13;	// <stdin>:5280:13
  wire [31:0] _T_14;	// <stdin>:5272:13
  wire [31:0] _T_15;	// <stdin>:5264:13
  wire [31:0] _T_16;	// <stdin>:5256:13
  wire [31:0] _T_17;	// <stdin>:5248:13
  wire [31:0] _T_18;	// <stdin>:5240:13
  wire [31:0] _T_19;	// <stdin>:5232:13
  wire [31:0] _T_20;	// <stdin>:5224:13
  wire [31:0] _T_21;	// <stdin>:5216:13
  wire [31:0] _T_22;	// <stdin>:5208:13
  wire [31:0] _T_23;	// <stdin>:5200:13
  wire [31:0] _T_24;	// <stdin>:5192:13
  wire [31:0] _T_25;	// <stdin>:5184:13
  wire [31:0] _T_26;	// <stdin>:5176:13
  wire [31:0] _T_27;	// <stdin>:5168:13
  wire [31:0] _T_28;	// <stdin>:5160:13
  wire [31:0] _T_29;	// <stdin>:5152:13
  wire [31:0] _T_30;	// <stdin>:5144:13
  wire [31:0] _T_31;	// <stdin>:5136:13
  wire [31:0] _T_32;	// <stdin>:5128:13
  wire [31:0] _T_33;	// <stdin>:5120:13
  wire [31:0] _T_34;	// <stdin>:5112:13
  wire [31:0] _T_35;	// <stdin>:5104:13
  wire [31:0] _T_36;	// <stdin>:5096:13
  wire [31:0] _T_37;	// <stdin>:5088:13
  wire [31:0] _T_38;	// <stdin>:5080:13
  wire [31:0] _T_39;	// <stdin>:5072:13
  wire [31:0] _T_40;	// <stdin>:5064:13
  wire [31:0] _T_41;	// <stdin>:5056:13
  wire [31:0] _T_42;	// <stdin>:5048:13
  wire [31:0] _T_43;	// <stdin>:5040:13
  wire [31:0] _T_44;	// <stdin>:5032:13
  wire [31:0] _T_45;	// <stdin>:5024:13
  wire [31:0] _T_46;	// <stdin>:5016:13
  wire [31:0] _T_47;	// <stdin>:5008:13
  wire [31:0] _T_48;	// <stdin>:5000:13
  wire [31:0] _T_49;	// <stdin>:4992:13
  wire [31:0] _T_50;	// <stdin>:4984:13
  wire [31:0] _T_51;	// <stdin>:4976:13
  wire [31:0] _T_52;	// <stdin>:4968:13
  wire [31:0] _T_53;	// <stdin>:4960:13
  wire [31:0] _T_54;	// <stdin>:4952:13
  wire [31:0] _T_55;	// <stdin>:4944:13
  wire [31:0] _T_56;	// <stdin>:4936:13
  wire [31:0] _T_57;	// <stdin>:4928:13
  wire [31:0] _T_58;	// <stdin>:4920:13
  wire [31:0] _T_59;	// <stdin>:4912:13
  wire [31:0] _T_60;	// <stdin>:4904:13
  wire [31:0] _T_61;	// <stdin>:4896:13
  wire [31:0] _T_62;	// <stdin>:4888:13
  wire [31:0] _T_63;	// <stdin>:4880:13
  wire [31:0] _T_64;	// <stdin>:4872:13
  wire [31:0] _T_65;	// <stdin>:4864:13
  wire [31:0] _T_66;	// <stdin>:4856:13
  wire [31:0] _T_67;	// <stdin>:4848:13
  wire [31:0] _T_68;	// <stdin>:4840:13
  wire [31:0] _T_69;	// <stdin>:4832:13
  wire [31:0] _T_70;	// <stdin>:4824:13
  wire [31:0] _T_71;	// <stdin>:4816:13
  wire [31:0] _T_72;	// <stdin>:4808:13
  wire [31:0] _T_73;	// <stdin>:4800:13
  wire [31:0] _T_74;	// <stdin>:4792:13
  wire [31:0] _T_75;	// <stdin>:4784:13
  wire [31:0] _T_76;	// <stdin>:4776:13
  wire [31:0] _T_77;	// <stdin>:4768:13
  wire [31:0] _T_78;	// <stdin>:4760:13
  wire [31:0] _T_79;	// <stdin>:4752:13
  wire [31:0] _T_80;	// <stdin>:4744:13
  wire [31:0] _T_81;	// <stdin>:4736:13
  wire [31:0] _T_82;	// <stdin>:4728:13
  wire [31:0] _T_83;	// <stdin>:4720:13
  wire [31:0] _T_84;	// <stdin>:4712:13
  wire [31:0] _T_85;	// <stdin>:4704:13
  wire [31:0] _T_86;	// <stdin>:4696:13
  wire [31:0] _T_87;	// <stdin>:4688:13
  wire [31:0] _T_88;	// <stdin>:4680:13
  wire [31:0] _T_89;	// <stdin>:4672:13
  wire [31:0] _T_90;	// <stdin>:4664:13
  wire [31:0] _T_91;	// <stdin>:4656:13
  wire [31:0] _T_92;	// <stdin>:4648:13
  wire [31:0] _T_93;	// <stdin>:4640:13
  wire [31:0] _T_94;	// <stdin>:4632:13
  wire [31:0] _T_95;	// <stdin>:4624:13
  wire [31:0] _T_96;	// <stdin>:4616:13
  wire [31:0] _T_97;	// <stdin>:4608:13
  wire [31:0] _T_98;	// <stdin>:4600:13
  wire [31:0] _T_99;	// <stdin>:4592:13
  wire [31:0] _T_100;	// <stdin>:4584:13
  wire [31:0] _T_101;	// <stdin>:4576:13
  wire [31:0] _T_102;	// <stdin>:4568:13
  wire [31:0] _T_103;	// <stdin>:4560:13
  wire [31:0] _T_104;	// <stdin>:4552:13
  wire [31:0] _T_105;	// <stdin>:4544:13
  wire [31:0] _T_106;	// <stdin>:4536:13
  wire [31:0] _T_107;	// <stdin>:4528:13
  wire [31:0] _T_108;	// <stdin>:4520:13
  wire [31:0] _T_109;	// <stdin>:4512:13
  wire [31:0] _T_110;	// <stdin>:4504:13
  wire [31:0] _T_111;	// <stdin>:4496:13
  wire [31:0] _T_112;	// <stdin>:4488:13
  wire [31:0] _T_113;	// <stdin>:4480:12
  wire [31:0] _T_114;	// <stdin>:4472:12
  wire [31:0] _T_115;	// <stdin>:4464:12
  wire [31:0] _T_116;	// <stdin>:4456:12
  wire [31:0] _T_117;	// <stdin>:4448:12
  wire [31:0] _T_118;	// <stdin>:4440:12
  wire [31:0] _T_119;	// <stdin>:4432:12
  wire [31:0] _T_120;	// <stdin>:4424:12
  wire [31:0] _T_121;	// <stdin>:4416:12
  wire [31:0] _T_122;	// <stdin>:4408:12
  wire [31:0] _T_123;	// <stdin>:4400:12
  wire [31:0] _T_124;	// <stdin>:4392:12
  wire [31:0] _T_125;	// <stdin>:4384:12
  wire [31:0] _T_126;	// <stdin>:4376:12
  wire [31:0] _T_127;	// <stdin>:4368:12
  wire [31:0] _T_128;	// <stdin>:4360:12
  wire [31:0] _T_129;	// <stdin>:4352:12
  wire [31:0] _T_130;	// <stdin>:4344:12
  wire [31:0] _T_131;	// <stdin>:4336:12
  wire [31:0] _T_132;	// <stdin>:4328:12
  wire [31:0] _T_133;	// <stdin>:4320:12
  wire [31:0] _T_134;	// <stdin>:4312:12
  wire [31:0] _T_135;	// <stdin>:4304:12
  wire [31:0] _T_136;	// <stdin>:4296:12
  wire [31:0] _T_137;	// <stdin>:4288:12
  wire [31:0] _T_138;	// <stdin>:4280:12
  wire [31:0] _T_139;	// <stdin>:4272:12
  wire [31:0] _T_140;	// <stdin>:4264:12
  wire [31:0] _T_141;	// <stdin>:4256:12
  wire [31:0] _T_142;	// <stdin>:4248:12
  wire [31:0] _T_143;	// <stdin>:4240:12
  wire [31:0] _T_144;	// <stdin>:4232:12
  wire [31:0] _T_145;	// <stdin>:4224:12
  wire [31:0] _T_146;	// <stdin>:4216:12
  wire [31:0] _T_147;	// <stdin>:4208:12
  wire [31:0] _T_148;	// <stdin>:4200:12
  wire [31:0] _T_149;	// <stdin>:4192:12
  wire [31:0] _T_150;	// <stdin>:4184:12
  wire [31:0] _T_151;	// <stdin>:4176:12
  wire [31:0] _T_152;	// <stdin>:4168:12
  wire [31:0] _T_153;	// <stdin>:4160:12
  wire [31:0] _T_154;	// <stdin>:4152:12
  wire [31:0] _T_155;	// <stdin>:4144:12
  wire [31:0] _T_156;	// <stdin>:4136:12
  wire [31:0] _T_157;	// <stdin>:4128:12
  wire [31:0] _T_158;	// <stdin>:4120:12
  wire [31:0] _T_159;	// <stdin>:4112:12
  wire [31:0] _T_160;	// <stdin>:4104:12
  wire [31:0] _T_161;	// <stdin>:4096:12
  wire [31:0] _T_162;	// <stdin>:4088:12
  wire [31:0] _T_163;	// <stdin>:4080:12
  wire [31:0] _T_164;	// <stdin>:4072:12
  wire [31:0] _T_165;	// <stdin>:4064:12
  wire [31:0] _T_166;	// <stdin>:4056:12
  wire [31:0] _T_167;	// <stdin>:4048:12
  wire [31:0] _T_168;	// <stdin>:4040:12
  wire [31:0] _T_169;	// <stdin>:4032:12
  wire [31:0] _T_170;	// <stdin>:4024:12
  wire [31:0] _T_171;	// <stdin>:4016:12
  wire [31:0] _T_172;	// <stdin>:4008:12
  wire [31:0] _T_173;	// <stdin>:4000:12
  wire [31:0] _T_174;	// <stdin>:3992:12
  wire [31:0] _T_175;	// <stdin>:3984:12
  wire [31:0] _T_176;	// <stdin>:3976:12
  wire [31:0] _T_177;	// <stdin>:3968:12
  wire [31:0] _T_178;	// <stdin>:3960:12
  wire [31:0] _T_179;	// <stdin>:3952:12
  wire [31:0] _T_180;	// <stdin>:3944:12
  wire [31:0] _T_181;	// <stdin>:3936:12
  wire [31:0] _T_182;	// <stdin>:3928:12
  wire [31:0] _T_183;	// <stdin>:3920:12
  wire [31:0] _T_184;	// <stdin>:3912:12
  wire [31:0] _T_185;	// <stdin>:3904:12
  wire [31:0] _T_186;	// <stdin>:3896:12
  wire [31:0] _T_187;	// <stdin>:3888:12
  wire [31:0] _T_188;	// <stdin>:3880:12
  wire [31:0] _T_189;	// <stdin>:3872:12
  wire [31:0] _T_190;	// <stdin>:3864:12
  wire [31:0] _T_191;	// <stdin>:3856:12
  wire [31:0] _T_192;	// <stdin>:3848:12
  wire [31:0] _T_193;	// <stdin>:3840:12
  wire [31:0] _T_194;	// <stdin>:3832:12
  wire [31:0] _T_195;	// <stdin>:3824:12
  wire [31:0] _T_196;	// <stdin>:3816:12
  wire [31:0] _T_197;	// <stdin>:3808:12
  wire [31:0] _T_198;	// <stdin>:3800:12
  wire [31:0] _T_199;	// <stdin>:3792:12
  wire [31:0] _T_200;	// <stdin>:3784:12
  wire [31:0] _T_201;	// <stdin>:3776:12
  wire [31:0] _T_202;	// <stdin>:3768:12
  wire [31:0] _T_203;	// <stdin>:3760:12
  wire [31:0] _T_204;	// <stdin>:3752:12
  wire [31:0] _T_205;	// <stdin>:3744:12
  wire [31:0] _T_206;	// <stdin>:3736:12
  wire [31:0] _T_207;	// <stdin>:3728:12
  wire [31:0] _T_208;	// <stdin>:3720:12
  wire [31:0] _T_209;	// <stdin>:3712:12
  wire [31:0] _T_210;	// <stdin>:3704:12
  wire [31:0] _T_211;	// <stdin>:3696:12
  wire [31:0] _T_212;	// <stdin>:3688:12
  wire [31:0] _T_213;	// <stdin>:3680:12
  wire [31:0] _T_214;	// <stdin>:3672:12
  wire [31:0] _T_215;	// <stdin>:3664:12
  wire [31:0] _T_216;	// <stdin>:3656:12
  wire [31:0] _T_217;	// <stdin>:3648:12
  wire [31:0] _T_218;	// <stdin>:3640:12
  wire [31:0] _T_219;	// <stdin>:3632:12
  wire [31:0] _T_220;	// <stdin>:3624:12
  wire [31:0] _T_221;	// <stdin>:3616:12
  wire [31:0] _T_222;	// <stdin>:3608:12
  wire [31:0] _T_223;	// <stdin>:3600:12
  wire [31:0] _T_224;	// <stdin>:3592:12
  wire [31:0] _T_225;	// <stdin>:3584:12
  wire [31:0] _T_226;	// <stdin>:3576:12
  wire [31:0] _T_227;	// <stdin>:3568:12
  wire [31:0] _T_228;	// <stdin>:3560:12
  wire [31:0] _T_229;	// <stdin>:3552:12
  wire [31:0] _T_230;	// <stdin>:3544:12
  wire [31:0] _T_231;	// <stdin>:3536:12
  wire [31:0] _T_232;	// <stdin>:3528:12
  wire [31:0] _T_233;	// <stdin>:3520:12
  wire [31:0] _T_234;	// <stdin>:3512:12
  wire [31:0] _T_235;	// <stdin>:3504:12
  wire [31:0] _T_236;	// <stdin>:3496:12
  wire [31:0] _T_237;	// <stdin>:3488:12
  wire [31:0] _T_238;	// <stdin>:3480:12
  wire [31:0] _T_239;	// <stdin>:3472:12
  wire [31:0] _T_240;	// <stdin>:3464:12
  wire [31:0] _T_241;	// <stdin>:3456:11
  wire [31:0] _T_242;	// <stdin>:3448:11
  wire [31:0] _T_243;	// <stdin>:3440:11
  wire [31:0] _T_244;	// <stdin>:3432:11
  wire [31:0] _T_245;	// <stdin>:3424:11
  wire [31:0] _T_246;	// <stdin>:3416:11
  wire [31:0] _T_247;	// <stdin>:3408:11
  wire [31:0] _T_248;	// <stdin>:3400:11
  wire [31:0] _T_249;	// <stdin>:3392:11
  wire [31:0] _T_250;	// <stdin>:3384:11
  wire [31:0] _T_251;	// <stdin>:3376:11
  wire [31:0] _T_252;	// <stdin>:3368:11
  wire [31:0] _T_253;	// <stdin>:3360:11
  wire [31:0] _T_254;	// <stdin>:3352:10
  reg  [31:0] Register_inst0;	// <stdin>:3351:23
  reg  [31:0] Register_inst1;	// <stdin>:3359:23
  reg  [31:0] Register_inst2;	// <stdin>:3367:23
  reg  [31:0] Register_inst3;	// <stdin>:3375:23
  reg  [31:0] Register_inst4;	// <stdin>:3383:23
  reg  [31:0] Register_inst5;	// <stdin>:3391:23
  reg  [31:0] Register_inst6;	// <stdin>:3399:23
  reg  [31:0] Register_inst7;	// <stdin>:3407:23
  reg  [31:0] Register_inst8;	// <stdin>:3415:23
  reg  [31:0] Register_inst9;	// <stdin>:3423:23
  reg  [31:0] Register_inst10;	// <stdin>:3431:24
  reg  [31:0] Register_inst11;	// <stdin>:3439:24
  reg  [31:0] Register_inst12;	// <stdin>:3447:24
  reg  [31:0] Register_inst13;	// <stdin>:3455:24
  reg  [31:0] Register_inst14;	// <stdin>:3463:24
  reg  [31:0] Register_inst15;	// <stdin>:3471:24
  reg  [31:0] Register_inst16;	// <stdin>:3479:24
  reg  [31:0] Register_inst17;	// <stdin>:3487:24
  reg  [31:0] Register_inst18;	// <stdin>:3495:24
  reg  [31:0] Register_inst19;	// <stdin>:3503:24
  reg  [31:0] Register_inst20;	// <stdin>:3511:24
  reg  [31:0] Register_inst21;	// <stdin>:3519:24
  reg  [31:0] Register_inst22;	// <stdin>:3527:24
  reg  [31:0] Register_inst23;	// <stdin>:3535:24
  reg  [31:0] Register_inst24;	// <stdin>:3543:24
  reg  [31:0] Register_inst25;	// <stdin>:3551:24
  reg  [31:0] Register_inst26;	// <stdin>:3559:24
  reg  [31:0] Register_inst27;	// <stdin>:3567:24
  reg  [31:0] Register_inst28;	// <stdin>:3575:24
  reg  [31:0] Register_inst29;	// <stdin>:3583:24
  reg  [31:0] Register_inst30;	// <stdin>:3591:24
  reg  [31:0] Register_inst31;	// <stdin>:3599:24
  reg  [31:0] Register_inst32;	// <stdin>:3607:24
  reg  [31:0] Register_inst33;	// <stdin>:3615:24
  reg  [31:0] Register_inst34;	// <stdin>:3623:24
  reg  [31:0] Register_inst35;	// <stdin>:3631:24
  reg  [31:0] Register_inst36;	// <stdin>:3639:24
  reg  [31:0] Register_inst37;	// <stdin>:3647:24
  reg  [31:0] Register_inst38;	// <stdin>:3655:24
  reg  [31:0] Register_inst39;	// <stdin>:3663:24
  reg  [31:0] Register_inst40;	// <stdin>:3671:24
  reg  [31:0] Register_inst41;	// <stdin>:3679:24
  reg  [31:0] Register_inst42;	// <stdin>:3687:24
  reg  [31:0] Register_inst43;	// <stdin>:3695:24
  reg  [31:0] Register_inst44;	// <stdin>:3703:24
  reg  [31:0] Register_inst45;	// <stdin>:3711:24
  reg  [31:0] Register_inst46;	// <stdin>:3719:24
  reg  [31:0] Register_inst47;	// <stdin>:3727:24
  reg  [31:0] Register_inst48;	// <stdin>:3735:24
  reg  [31:0] Register_inst49;	// <stdin>:3743:24
  reg  [31:0] Register_inst50;	// <stdin>:3751:24
  reg  [31:0] Register_inst51;	// <stdin>:3759:24
  reg  [31:0] Register_inst52;	// <stdin>:3767:24
  reg  [31:0] Register_inst53;	// <stdin>:3775:24
  reg  [31:0] Register_inst54;	// <stdin>:3783:24
  reg  [31:0] Register_inst55;	// <stdin>:3791:24
  reg  [31:0] Register_inst56;	// <stdin>:3799:24
  reg  [31:0] Register_inst57;	// <stdin>:3807:24
  reg  [31:0] Register_inst58;	// <stdin>:3815:24
  reg  [31:0] Register_inst59;	// <stdin>:3823:24
  reg  [31:0] Register_inst60;	// <stdin>:3831:24
  reg  [31:0] Register_inst61;	// <stdin>:3839:24
  reg  [31:0] Register_inst62;	// <stdin>:3847:24
  reg  [31:0] Register_inst63;	// <stdin>:3855:24
  reg  [31:0] Register_inst64;	// <stdin>:3863:24
  reg  [31:0] Register_inst65;	// <stdin>:3871:24
  reg  [31:0] Register_inst66;	// <stdin>:3879:24
  reg  [31:0] Register_inst67;	// <stdin>:3887:24
  reg  [31:0] Register_inst68;	// <stdin>:3895:24
  reg  [31:0] Register_inst69;	// <stdin>:3903:24
  reg  [31:0] Register_inst70;	// <stdin>:3911:24
  reg  [31:0] Register_inst71;	// <stdin>:3919:24
  reg  [31:0] Register_inst72;	// <stdin>:3927:24
  reg  [31:0] Register_inst73;	// <stdin>:3935:24
  reg  [31:0] Register_inst74;	// <stdin>:3943:24
  reg  [31:0] Register_inst75;	// <stdin>:3951:24
  reg  [31:0] Register_inst76;	// <stdin>:3959:24
  reg  [31:0] Register_inst77;	// <stdin>:3967:24
  reg  [31:0] Register_inst78;	// <stdin>:3975:24
  reg  [31:0] Register_inst79;	// <stdin>:3983:24
  reg  [31:0] Register_inst80;	// <stdin>:3991:24
  reg  [31:0] Register_inst81;	// <stdin>:3999:24
  reg  [31:0] Register_inst82;	// <stdin>:4007:24
  reg  [31:0] Register_inst83;	// <stdin>:4015:24
  reg  [31:0] Register_inst84;	// <stdin>:4023:24
  reg  [31:0] Register_inst85;	// <stdin>:4031:24
  reg  [31:0] Register_inst86;	// <stdin>:4039:24
  reg  [31:0] Register_inst87;	// <stdin>:4047:24
  reg  [31:0] Register_inst88;	// <stdin>:4055:24
  reg  [31:0] Register_inst89;	// <stdin>:4063:24
  reg  [31:0] Register_inst90;	// <stdin>:4071:24
  reg  [31:0] Register_inst91;	// <stdin>:4079:24
  reg  [31:0] Register_inst92;	// <stdin>:4087:24
  reg  [31:0] Register_inst93;	// <stdin>:4095:24
  reg  [31:0] Register_inst94;	// <stdin>:4103:24
  reg  [31:0] Register_inst95;	// <stdin>:4111:24
  reg  [31:0] Register_inst96;	// <stdin>:4119:24
  reg  [31:0] Register_inst97;	// <stdin>:4127:24
  reg  [31:0] Register_inst98;	// <stdin>:4135:24
  reg  [31:0] Register_inst99;	// <stdin>:4143:24
  reg  [31:0] Register_inst100;	// <stdin>:4151:25
  reg  [31:0] Register_inst101;	// <stdin>:4159:25
  reg  [31:0] Register_inst102;	// <stdin>:4167:25
  reg  [31:0] Register_inst103;	// <stdin>:4175:25
  reg  [31:0] Register_inst104;	// <stdin>:4183:25
  reg  [31:0] Register_inst105;	// <stdin>:4191:25
  reg  [31:0] Register_inst106;	// <stdin>:4199:25
  reg  [31:0] Register_inst107;	// <stdin>:4207:25
  reg  [31:0] Register_inst108;	// <stdin>:4215:25
  reg  [31:0] Register_inst109;	// <stdin>:4223:25
  reg  [31:0] Register_inst110;	// <stdin>:4231:25
  reg  [31:0] Register_inst111;	// <stdin>:4239:25
  reg  [31:0] Register_inst112;	// <stdin>:4247:25
  reg  [31:0] Register_inst113;	// <stdin>:4255:25
  reg  [31:0] Register_inst114;	// <stdin>:4263:25
  reg  [31:0] Register_inst115;	// <stdin>:4271:25
  reg  [31:0] Register_inst116;	// <stdin>:4279:25
  reg  [31:0] Register_inst117;	// <stdin>:4287:25
  reg  [31:0] Register_inst118;	// <stdin>:4295:25
  reg  [31:0] Register_inst119;	// <stdin>:4303:25
  reg  [31:0] Register_inst120;	// <stdin>:4311:25
  reg  [31:0] Register_inst121;	// <stdin>:4319:25
  reg  [31:0] Register_inst122;	// <stdin>:4327:25
  reg  [31:0] Register_inst123;	// <stdin>:4335:25
  reg  [31:0] Register_inst124;	// <stdin>:4343:25
  reg  [31:0] Register_inst125;	// <stdin>:4351:25
  reg  [31:0] Register_inst126;	// <stdin>:4359:25
  reg  [31:0] Register_inst127;	// <stdin>:4367:25
  reg  [31:0] Register_inst128;	// <stdin>:4375:25
  reg  [31:0] Register_inst129;	// <stdin>:4383:25
  reg  [31:0] Register_inst130;	// <stdin>:4391:25
  reg  [31:0] Register_inst131;	// <stdin>:4399:25
  reg  [31:0] Register_inst132;	// <stdin>:4407:25
  reg  [31:0] Register_inst133;	// <stdin>:4415:25
  reg  [31:0] Register_inst134;	// <stdin>:4423:25
  reg  [31:0] Register_inst135;	// <stdin>:4431:25
  reg  [31:0] Register_inst136;	// <stdin>:4439:25
  reg  [31:0] Register_inst137;	// <stdin>:4447:25
  reg  [31:0] Register_inst138;	// <stdin>:4455:25
  reg  [31:0] Register_inst139;	// <stdin>:4463:25
  reg  [31:0] Register_inst140;	// <stdin>:4471:25
  reg  [31:0] Register_inst141;	// <stdin>:4479:25
  reg  [31:0] Register_inst142;	// <stdin>:4487:25
  reg  [31:0] Register_inst143;	// <stdin>:4495:25
  reg  [31:0] Register_inst144;	// <stdin>:4503:25
  reg  [31:0] Register_inst145;	// <stdin>:4511:25
  reg  [31:0] Register_inst146;	// <stdin>:4519:25
  reg  [31:0] Register_inst147;	// <stdin>:4527:25
  reg  [31:0] Register_inst148;	// <stdin>:4535:25
  reg  [31:0] Register_inst149;	// <stdin>:4543:25
  reg  [31:0] Register_inst150;	// <stdin>:4551:25
  reg  [31:0] Register_inst151;	// <stdin>:4559:25
  reg  [31:0] Register_inst152;	// <stdin>:4567:25
  reg  [31:0] Register_inst153;	// <stdin>:4575:25
  reg  [31:0] Register_inst154;	// <stdin>:4583:25
  reg  [31:0] Register_inst155;	// <stdin>:4591:25
  reg  [31:0] Register_inst156;	// <stdin>:4599:25
  reg  [31:0] Register_inst157;	// <stdin>:4607:25
  reg  [31:0] Register_inst158;	// <stdin>:4615:25
  reg  [31:0] Register_inst159;	// <stdin>:4623:25
  reg  [31:0] Register_inst160;	// <stdin>:4631:25
  reg  [31:0] Register_inst161;	// <stdin>:4639:25
  reg  [31:0] Register_inst162;	// <stdin>:4647:25
  reg  [31:0] Register_inst163;	// <stdin>:4655:25
  reg  [31:0] Register_inst164;	// <stdin>:4663:25
  reg  [31:0] Register_inst165;	// <stdin>:4671:25
  reg  [31:0] Register_inst166;	// <stdin>:4679:25
  reg  [31:0] Register_inst167;	// <stdin>:4687:25
  reg  [31:0] Register_inst168;	// <stdin>:4695:25
  reg  [31:0] Register_inst169;	// <stdin>:4703:25
  reg  [31:0] Register_inst170;	// <stdin>:4711:25
  reg  [31:0] Register_inst171;	// <stdin>:4719:25
  reg  [31:0] Register_inst172;	// <stdin>:4727:25
  reg  [31:0] Register_inst173;	// <stdin>:4735:25
  reg  [31:0] Register_inst174;	// <stdin>:4743:25
  reg  [31:0] Register_inst175;	// <stdin>:4751:25
  reg  [31:0] Register_inst176;	// <stdin>:4759:25
  reg  [31:0] Register_inst177;	// <stdin>:4767:25
  reg  [31:0] Register_inst178;	// <stdin>:4775:25
  reg  [31:0] Register_inst179;	// <stdin>:4783:25
  reg  [31:0] Register_inst180;	// <stdin>:4791:25
  reg  [31:0] Register_inst181;	// <stdin>:4799:25
  reg  [31:0] Register_inst182;	// <stdin>:4807:25
  reg  [31:0] Register_inst183;	// <stdin>:4815:25
  reg  [31:0] Register_inst184;	// <stdin>:4823:25
  reg  [31:0] Register_inst185;	// <stdin>:4831:25
  reg  [31:0] Register_inst186;	// <stdin>:4839:25
  reg  [31:0] Register_inst187;	// <stdin>:4847:25
  reg  [31:0] Register_inst188;	// <stdin>:4855:25
  reg  [31:0] Register_inst189;	// <stdin>:4863:25
  reg  [31:0] Register_inst190;	// <stdin>:4871:25
  reg  [31:0] Register_inst191;	// <stdin>:4879:25
  reg  [31:0] Register_inst192;	// <stdin>:4887:25
  reg  [31:0] Register_inst193;	// <stdin>:4895:25
  reg  [31:0] Register_inst194;	// <stdin>:4903:25
  reg  [31:0] Register_inst195;	// <stdin>:4911:25
  reg  [31:0] Register_inst196;	// <stdin>:4919:25
  reg  [31:0] Register_inst197;	// <stdin>:4927:25
  reg  [31:0] Register_inst198;	// <stdin>:4935:25
  reg  [31:0] Register_inst199;	// <stdin>:4943:25
  reg  [31:0] Register_inst200;	// <stdin>:4951:25
  reg  [31:0] Register_inst201;	// <stdin>:4959:25
  reg  [31:0] Register_inst202;	// <stdin>:4967:25
  reg  [31:0] Register_inst203;	// <stdin>:4975:25
  reg  [31:0] Register_inst204;	// <stdin>:4983:25
  reg  [31:0] Register_inst205;	// <stdin>:4991:25
  reg  [31:0] Register_inst206;	// <stdin>:4999:25
  reg  [31:0] Register_inst207;	// <stdin>:5007:25
  reg  [31:0] Register_inst208;	// <stdin>:5015:25
  reg  [31:0] Register_inst209;	// <stdin>:5023:25
  reg  [31:0] Register_inst210;	// <stdin>:5031:25
  reg  [31:0] Register_inst211;	// <stdin>:5039:25
  reg  [31:0] Register_inst212;	// <stdin>:5047:25
  reg  [31:0] Register_inst213;	// <stdin>:5055:25
  reg  [31:0] Register_inst214;	// <stdin>:5063:25
  reg  [31:0] Register_inst215;	// <stdin>:5071:25
  reg  [31:0] Register_inst216;	// <stdin>:5079:25
  reg  [31:0] Register_inst217;	// <stdin>:5087:25
  reg  [31:0] Register_inst218;	// <stdin>:5095:25
  reg  [31:0] Register_inst219;	// <stdin>:5103:25
  reg  [31:0] Register_inst220;	// <stdin>:5111:25
  reg  [31:0] Register_inst221;	// <stdin>:5119:25
  reg  [31:0] Register_inst222;	// <stdin>:5127:25
  reg  [31:0] Register_inst223;	// <stdin>:5135:25
  reg  [31:0] Register_inst224;	// <stdin>:5143:25
  reg  [31:0] Register_inst225;	// <stdin>:5151:25
  reg  [31:0] Register_inst226;	// <stdin>:5159:25
  reg  [31:0] Register_inst227;	// <stdin>:5167:25
  reg  [31:0] Register_inst228;	// <stdin>:5175:25
  reg  [31:0] Register_inst229;	// <stdin>:5183:25
  reg  [31:0] Register_inst230;	// <stdin>:5191:25
  reg  [31:0] Register_inst231;	// <stdin>:5199:25
  reg  [31:0] Register_inst232;	// <stdin>:5207:25
  reg  [31:0] Register_inst233;	// <stdin>:5215:25
  reg  [31:0] Register_inst234;	// <stdin>:5223:25
  reg  [31:0] Register_inst235;	// <stdin>:5231:25
  reg  [31:0] Register_inst236;	// <stdin>:5239:25
  reg  [31:0] Register_inst237;	// <stdin>:5247:25
  reg  [31:0] Register_inst238;	// <stdin>:5255:25
  reg  [31:0] Register_inst239;	// <stdin>:5263:25
  reg  [31:0] Register_inst240;	// <stdin>:5271:25
  reg  [31:0] Register_inst241;	// <stdin>:5279:25
  reg  [31:0] Register_inst242;	// <stdin>:5287:25
  reg  [31:0] Register_inst243;	// <stdin>:5295:25
  reg  [31:0] Register_inst244;	// <stdin>:5303:25
  reg  [31:0] Register_inst245;	// <stdin>:5311:25
  reg  [31:0] Register_inst246;	// <stdin>:5319:25
  reg  [31:0] Register_inst247;	// <stdin>:5327:25
  reg  [31:0] Register_inst248;	// <stdin>:5335:25
  reg  [31:0] Register_inst249;	// <stdin>:5343:25
  reg  [31:0] Register_inst250;	// <stdin>:5351:25
  reg  [31:0] Register_inst251;	// <stdin>:5359:25
  reg  [31:0] Register_inst252;	// <stdin>:5367:25
  reg  [31:0] Register_inst253;	// <stdin>:5375:25
  reg  [31:0] Register_inst254;	// <stdin>:5383:25
  reg  [31:0] Register_inst255;	// <stdin>:5391:25

  wire [31:0] _T_255 = ({{_T_254}, {write_0.data}})[write_0.addr == 8'h0 & write_0_en];	// <stdin>:3344:14, :3345:10, :3346:10, :3347:10, :3348:10, :3349:10, :3350:10, :3352:10
  assign _T_254 = Register_inst0;	// <stdin>:3352:10
  wire [31:0] _T_256 = ({{_T_253}, {write_0.data}})[write_0.addr == 8'h1 & write_0_en];	// <stdin>:3343:14, :3353:10, :3354:10, :3355:10, :3356:11, :3357:11, :3358:11, :3360:11
  assign _T_253 = Register_inst1;	// <stdin>:3360:11
  wire [31:0] _T_257 = ({{_T_252}, {write_0.data}})[write_0.addr == 8'h2 & write_0_en];	// <stdin>:3342:14, :3361:11, :3362:11, :3363:11, :3364:11, :3365:11, :3366:11, :3368:11
  assign _T_252 = Register_inst2;	// <stdin>:3368:11
  wire [31:0] _T_258 = ({{_T_251}, {write_0.data}})[write_0.addr == 8'h3 & write_0_en];	// <stdin>:3341:14, :3369:11, :3370:11, :3371:11, :3372:11, :3373:11, :3374:11, :3376:11
  assign _T_251 = Register_inst3;	// <stdin>:3376:11
  wire [31:0] _T_259 = ({{_T_250}, {write_0.data}})[write_0.addr == 8'h4 & write_0_en];	// <stdin>:3340:14, :3377:11, :3378:11, :3379:11, :3380:11, :3381:11, :3382:11, :3384:11
  assign _T_250 = Register_inst4;	// <stdin>:3384:11
  wire [31:0] _T_260 = ({{_T_249}, {write_0.data}})[write_0.addr == 8'h5 & write_0_en];	// <stdin>:3339:14, :3385:11, :3386:11, :3387:11, :3388:11, :3389:11, :3390:11, :3392:11
  assign _T_249 = Register_inst5;	// <stdin>:3392:11
  wire [31:0] _T_261 = ({{_T_248}, {write_0.data}})[write_0.addr == 8'h6 & write_0_en];	// <stdin>:3338:14, :3393:11, :3394:11, :3395:11, :3396:11, :3397:11, :3398:11, :3400:11
  assign _T_248 = Register_inst6;	// <stdin>:3400:11
  wire [31:0] _T_262 = ({{_T_247}, {write_0.data}})[write_0.addr == 8'h7 & write_0_en];	// <stdin>:3337:14, :3401:11, :3402:11, :3403:11, :3404:11, :3405:11, :3406:11, :3408:11
  assign _T_247 = Register_inst7;	// <stdin>:3408:11
  wire [31:0] _T_263 = ({{_T_246}, {write_0.data}})[write_0.addr == 8'h8 & write_0_en];	// <stdin>:3336:14, :3409:11, :3410:11, :3411:11, :3412:11, :3413:11, :3414:11, :3416:11
  assign _T_246 = Register_inst8;	// <stdin>:3416:11
  wire [31:0] _T_264 = ({{_T_245}, {write_0.data}})[write_0.addr == 8'h9 & write_0_en];	// <stdin>:3335:14, :3417:11, :3418:11, :3419:11, :3420:11, :3421:11, :3422:11, :3424:11
  assign _T_245 = Register_inst9;	// <stdin>:3424:11
  wire [31:0] _T_265 = ({{_T_244}, {write_0.data}})[write_0.addr == 8'hA & write_0_en];	// <stdin>:3334:15, :3425:11, :3426:11, :3427:11, :3428:11, :3429:11, :3430:11, :3432:11
  assign _T_244 = Register_inst10;	// <stdin>:3432:11
  wire [31:0] _T_266 = ({{_T_243}, {write_0.data}})[write_0.addr == 8'hB & write_0_en];	// <stdin>:3333:15, :3433:11, :3434:11, :3435:11, :3436:11, :3437:11, :3438:11, :3440:11
  assign _T_243 = Register_inst11;	// <stdin>:3440:11
  wire [31:0] _T_267 = ({{_T_242}, {write_0.data}})[write_0.addr == 8'hC & write_0_en];	// <stdin>:3332:15, :3441:11, :3442:11, :3443:11, :3444:11, :3445:11, :3446:11, :3448:11
  assign _T_242 = Register_inst12;	// <stdin>:3448:11
  wire [31:0] _T_268 = ({{_T_241}, {write_0.data}})[write_0.addr == 8'hD & write_0_en];	// <stdin>:3331:15, :3449:11, :3450:11, :3451:11, :3452:11, :3453:11, :3454:11, :3456:11
  assign _T_241 = Register_inst13;	// <stdin>:3456:11
  wire [31:0] _T_269 = ({{_T_240}, {write_0.data}})[write_0.addr == 8'hE & write_0_en];	// <stdin>:3330:15, :3457:11, :3458:11, :3459:12, :3460:12, :3461:12, :3462:12, :3464:12
  assign _T_240 = Register_inst14;	// <stdin>:3464:12
  wire [31:0] _T_270 = ({{_T_239}, {write_0.data}})[write_0.addr == 8'hF & write_0_en];	// <stdin>:3329:15, :3465:12, :3466:12, :3467:12, :3468:12, :3469:12, :3470:12, :3472:12
  assign _T_239 = Register_inst15;	// <stdin>:3472:12
  wire [31:0] _T_271 = ({{_T_238}, {write_0.data}})[write_0.addr == 8'h10 & write_0_en];	// <stdin>:3328:15, :3473:12, :3474:12, :3475:12, :3476:12, :3477:12, :3478:12, :3480:12
  assign _T_238 = Register_inst16;	// <stdin>:3480:12
  wire [31:0] _T_272 = ({{_T_237}, {write_0.data}})[write_0.addr == 8'h11 & write_0_en];	// <stdin>:3327:15, :3481:12, :3482:12, :3483:12, :3484:12, :3485:12, :3486:12, :3488:12
  assign _T_237 = Register_inst17;	// <stdin>:3488:12
  wire [31:0] _T_273 = ({{_T_236}, {write_0.data}})[write_0.addr == 8'h12 & write_0_en];	// <stdin>:3326:15, :3489:12, :3490:12, :3491:12, :3492:12, :3493:12, :3494:12, :3496:12
  assign _T_236 = Register_inst18;	// <stdin>:3496:12
  wire [31:0] _T_274 = ({{_T_235}, {write_0.data}})[write_0.addr == 8'h13 & write_0_en];	// <stdin>:3325:15, :3497:12, :3498:12, :3499:12, :3500:12, :3501:12, :3502:12, :3504:12
  assign _T_235 = Register_inst19;	// <stdin>:3504:12
  wire [31:0] _T_275 = ({{_T_234}, {write_0.data}})[write_0.addr == 8'h14 & write_0_en];	// <stdin>:3324:15, :3505:12, :3506:12, :3507:12, :3508:12, :3509:12, :3510:12, :3512:12
  assign _T_234 = Register_inst20;	// <stdin>:3512:12
  wire [31:0] _T_276 = ({{_T_233}, {write_0.data}})[write_0.addr == 8'h15 & write_0_en];	// <stdin>:3323:15, :3513:12, :3514:12, :3515:12, :3516:12, :3517:12, :3518:12, :3520:12
  assign _T_233 = Register_inst21;	// <stdin>:3520:12
  wire [31:0] _T_277 = ({{_T_232}, {write_0.data}})[write_0.addr == 8'h16 & write_0_en];	// <stdin>:3322:15, :3521:12, :3522:12, :3523:12, :3524:12, :3525:12, :3526:12, :3528:12
  assign _T_232 = Register_inst22;	// <stdin>:3528:12
  wire [31:0] _T_278 = ({{_T_231}, {write_0.data}})[write_0.addr == 8'h17 & write_0_en];	// <stdin>:3321:15, :3529:12, :3530:12, :3531:12, :3532:12, :3533:12, :3534:12, :3536:12
  assign _T_231 = Register_inst23;	// <stdin>:3536:12
  wire [31:0] _T_279 = ({{_T_230}, {write_0.data}})[write_0.addr == 8'h18 & write_0_en];	// <stdin>:3320:15, :3537:12, :3538:12, :3539:12, :3540:12, :3541:12, :3542:12, :3544:12
  assign _T_230 = Register_inst24;	// <stdin>:3544:12
  wire [31:0] _T_280 = ({{_T_229}, {write_0.data}})[write_0.addr == 8'h19 & write_0_en];	// <stdin>:3319:15, :3545:12, :3546:12, :3547:12, :3548:12, :3549:12, :3550:12, :3552:12
  assign _T_229 = Register_inst25;	// <stdin>:3552:12
  wire [31:0] _T_281 = ({{_T_228}, {write_0.data}})[write_0.addr == 8'h1A & write_0_en];	// <stdin>:3318:15, :3553:12, :3554:12, :3555:12, :3556:12, :3557:12, :3558:12, :3560:12
  assign _T_228 = Register_inst26;	// <stdin>:3560:12
  wire [31:0] _T_282 = ({{_T_227}, {write_0.data}})[write_0.addr == 8'h1B & write_0_en];	// <stdin>:3317:15, :3561:12, :3562:12, :3563:12, :3564:12, :3565:12, :3566:12, :3568:12
  assign _T_227 = Register_inst27;	// <stdin>:3568:12
  wire [31:0] _T_283 = ({{_T_226}, {write_0.data}})[write_0.addr == 8'h1C & write_0_en];	// <stdin>:3316:15, :3569:12, :3570:12, :3571:12, :3572:12, :3573:12, :3574:12, :3576:12
  assign _T_226 = Register_inst28;	// <stdin>:3576:12
  wire [31:0] _T_284 = ({{_T_225}, {write_0.data}})[write_0.addr == 8'h1D & write_0_en];	// <stdin>:3315:15, :3577:12, :3578:12, :3579:12, :3580:12, :3581:12, :3582:12, :3584:12
  assign _T_225 = Register_inst29;	// <stdin>:3584:12
  wire [31:0] _T_285 = ({{_T_224}, {write_0.data}})[write_0.addr == 8'h1E & write_0_en];	// <stdin>:3314:15, :3585:12, :3586:12, :3587:12, :3588:12, :3589:12, :3590:12, :3592:12
  assign _T_224 = Register_inst30;	// <stdin>:3592:12
  wire [31:0] _T_286 = ({{_T_223}, {write_0.data}})[write_0.addr == 8'h1F & write_0_en];	// <stdin>:3313:15, :3593:12, :3594:12, :3595:12, :3596:12, :3597:12, :3598:12, :3600:12
  assign _T_223 = Register_inst31;	// <stdin>:3600:12
  wire [31:0] _T_287 = ({{_T_222}, {write_0.data}})[write_0.addr == 8'h20 & write_0_en];	// <stdin>:3312:15, :3601:12, :3602:12, :3603:12, :3604:12, :3605:12, :3606:12, :3608:12
  assign _T_222 = Register_inst32;	// <stdin>:3608:12
  wire [31:0] _T_288 = ({{_T_221}, {write_0.data}})[write_0.addr == 8'h21 & write_0_en];	// <stdin>:3311:15, :3609:12, :3610:12, :3611:12, :3612:12, :3613:12, :3614:12, :3616:12
  assign _T_221 = Register_inst33;	// <stdin>:3616:12
  wire [31:0] _T_289 = ({{_T_220}, {write_0.data}})[write_0.addr == 8'h22 & write_0_en];	// <stdin>:3310:15, :3617:12, :3618:12, :3619:12, :3620:12, :3621:12, :3622:12, :3624:12
  assign _T_220 = Register_inst34;	// <stdin>:3624:12
  wire [31:0] _T_290 = ({{_T_219}, {write_0.data}})[write_0.addr == 8'h23 & write_0_en];	// <stdin>:3309:15, :3625:12, :3626:12, :3627:12, :3628:12, :3629:12, :3630:12, :3632:12
  assign _T_219 = Register_inst35;	// <stdin>:3632:12
  wire [31:0] _T_291 = ({{_T_218}, {write_0.data}})[write_0.addr == 8'h24 & write_0_en];	// <stdin>:3308:15, :3633:12, :3634:12, :3635:12, :3636:12, :3637:12, :3638:12, :3640:12
  assign _T_218 = Register_inst36;	// <stdin>:3640:12
  wire [31:0] _T_292 = ({{_T_217}, {write_0.data}})[write_0.addr == 8'h25 & write_0_en];	// <stdin>:3307:15, :3641:12, :3642:12, :3643:12, :3644:12, :3645:12, :3646:12, :3648:12
  assign _T_217 = Register_inst37;	// <stdin>:3648:12
  wire [31:0] _T_293 = ({{_T_216}, {write_0.data}})[write_0.addr == 8'h26 & write_0_en];	// <stdin>:3306:15, :3649:12, :3650:12, :3651:12, :3652:12, :3653:12, :3654:12, :3656:12
  assign _T_216 = Register_inst38;	// <stdin>:3656:12
  wire [31:0] _T_294 = ({{_T_215}, {write_0.data}})[write_0.addr == 8'h27 & write_0_en];	// <stdin>:3305:15, :3657:12, :3658:12, :3659:12, :3660:12, :3661:12, :3662:12, :3664:12
  assign _T_215 = Register_inst39;	// <stdin>:3664:12
  wire [31:0] _T_295 = ({{_T_214}, {write_0.data}})[write_0.addr == 8'h28 & write_0_en];	// <stdin>:3304:15, :3665:12, :3666:12, :3667:12, :3668:12, :3669:12, :3670:12, :3672:12
  assign _T_214 = Register_inst40;	// <stdin>:3672:12
  wire [31:0] _T_296 = ({{_T_213}, {write_0.data}})[write_0.addr == 8'h29 & write_0_en];	// <stdin>:3303:15, :3673:12, :3674:12, :3675:12, :3676:12, :3677:12, :3678:12, :3680:12
  assign _T_213 = Register_inst41;	// <stdin>:3680:12
  wire [31:0] _T_297 = ({{_T_212}, {write_0.data}})[write_0.addr == 8'h2A & write_0_en];	// <stdin>:3302:15, :3681:12, :3682:12, :3683:12, :3684:12, :3685:12, :3686:12, :3688:12
  assign _T_212 = Register_inst42;	// <stdin>:3688:12
  wire [31:0] _T_298 = ({{_T_211}, {write_0.data}})[write_0.addr == 8'h2B & write_0_en];	// <stdin>:3301:15, :3689:12, :3690:12, :3691:12, :3692:12, :3693:12, :3694:12, :3696:12
  assign _T_211 = Register_inst43;	// <stdin>:3696:12
  wire [31:0] _T_299 = ({{_T_210}, {write_0.data}})[write_0.addr == 8'h2C & write_0_en];	// <stdin>:3300:15, :3697:12, :3698:12, :3699:12, :3700:12, :3701:12, :3702:12, :3704:12
  assign _T_210 = Register_inst44;	// <stdin>:3704:12
  wire [31:0] _T_300 = ({{_T_209}, {write_0.data}})[write_0.addr == 8'h2D & write_0_en];	// <stdin>:3299:15, :3705:12, :3706:12, :3707:12, :3708:12, :3709:12, :3710:12, :3712:12
  assign _T_209 = Register_inst45;	// <stdin>:3712:12
  wire [31:0] _T_301 = ({{_T_208}, {write_0.data}})[write_0.addr == 8'h2E & write_0_en];	// <stdin>:3298:15, :3713:12, :3714:12, :3715:12, :3716:12, :3717:12, :3718:12, :3720:12
  assign _T_208 = Register_inst46;	// <stdin>:3720:12
  wire [31:0] _T_302 = ({{_T_207}, {write_0.data}})[write_0.addr == 8'h2F & write_0_en];	// <stdin>:3297:15, :3721:12, :3722:12, :3723:12, :3724:12, :3725:12, :3726:12, :3728:12
  assign _T_207 = Register_inst47;	// <stdin>:3728:12
  wire [31:0] _T_303 = ({{_T_206}, {write_0.data}})[write_0.addr == 8'h30 & write_0_en];	// <stdin>:3296:15, :3729:12, :3730:12, :3731:12, :3732:12, :3733:12, :3734:12, :3736:12
  assign _T_206 = Register_inst48;	// <stdin>:3736:12
  wire [31:0] _T_304 = ({{_T_205}, {write_0.data}})[write_0.addr == 8'h31 & write_0_en];	// <stdin>:3295:15, :3737:12, :3738:12, :3739:12, :3740:12, :3741:12, :3742:12, :3744:12
  assign _T_205 = Register_inst49;	// <stdin>:3744:12
  wire [31:0] _T_305 = ({{_T_204}, {write_0.data}})[write_0.addr == 8'h32 & write_0_en];	// <stdin>:3294:15, :3745:12, :3746:12, :3747:12, :3748:12, :3749:12, :3750:12, :3752:12
  assign _T_204 = Register_inst50;	// <stdin>:3752:12
  wire [31:0] _T_306 = ({{_T_203}, {write_0.data}})[write_0.addr == 8'h33 & write_0_en];	// <stdin>:3293:15, :3753:12, :3754:12, :3755:12, :3756:12, :3757:12, :3758:12, :3760:12
  assign _T_203 = Register_inst51;	// <stdin>:3760:12
  wire [31:0] _T_307 = ({{_T_202}, {write_0.data}})[write_0.addr == 8'h34 & write_0_en];	// <stdin>:3292:15, :3761:12, :3762:12, :3763:12, :3764:12, :3765:12, :3766:12, :3768:12
  assign _T_202 = Register_inst52;	// <stdin>:3768:12
  wire [31:0] _T_308 = ({{_T_201}, {write_0.data}})[write_0.addr == 8'h35 & write_0_en];	// <stdin>:3291:15, :3769:12, :3770:12, :3771:12, :3772:12, :3773:12, :3774:12, :3776:12
  assign _T_201 = Register_inst53;	// <stdin>:3776:12
  wire [31:0] _T_309 = ({{_T_200}, {write_0.data}})[write_0.addr == 8'h36 & write_0_en];	// <stdin>:3290:15, :3777:12, :3778:12, :3779:12, :3780:12, :3781:12, :3782:12, :3784:12
  assign _T_200 = Register_inst54;	// <stdin>:3784:12
  wire [31:0] _T_310 = ({{_T_199}, {write_0.data}})[write_0.addr == 8'h37 & write_0_en];	// <stdin>:3289:15, :3785:12, :3786:12, :3787:12, :3788:12, :3789:12, :3790:12, :3792:12
  assign _T_199 = Register_inst55;	// <stdin>:3792:12
  wire [31:0] _T_311 = ({{_T_198}, {write_0.data}})[write_0.addr == 8'h38 & write_0_en];	// <stdin>:3288:15, :3793:12, :3794:12, :3795:12, :3796:12, :3797:12, :3798:12, :3800:12
  assign _T_198 = Register_inst56;	// <stdin>:3800:12
  wire [31:0] _T_312 = ({{_T_197}, {write_0.data}})[write_0.addr == 8'h39 & write_0_en];	// <stdin>:3287:15, :3801:12, :3802:12, :3803:12, :3804:12, :3805:12, :3806:12, :3808:12
  assign _T_197 = Register_inst57;	// <stdin>:3808:12
  wire [31:0] _T_313 = ({{_T_196}, {write_0.data}})[write_0.addr == 8'h3A & write_0_en];	// <stdin>:3286:15, :3809:12, :3810:12, :3811:12, :3812:12, :3813:12, :3814:12, :3816:12
  assign _T_196 = Register_inst58;	// <stdin>:3816:12
  wire [31:0] _T_314 = ({{_T_195}, {write_0.data}})[write_0.addr == 8'h3B & write_0_en];	// <stdin>:3285:15, :3817:12, :3818:12, :3819:12, :3820:12, :3821:12, :3822:12, :3824:12
  assign _T_195 = Register_inst59;	// <stdin>:3824:12
  wire [31:0] _T_315 = ({{_T_194}, {write_0.data}})[write_0.addr == 8'h3C & write_0_en];	// <stdin>:3284:15, :3825:12, :3826:12, :3827:12, :3828:12, :3829:12, :3830:12, :3832:12
  assign _T_194 = Register_inst60;	// <stdin>:3832:12
  wire [31:0] _T_316 = ({{_T_193}, {write_0.data}})[write_0.addr == 8'h3D & write_0_en];	// <stdin>:3283:15, :3833:12, :3834:12, :3835:12, :3836:12, :3837:12, :3838:12, :3840:12
  assign _T_193 = Register_inst61;	// <stdin>:3840:12
  wire [31:0] _T_317 = ({{_T_192}, {write_0.data}})[write_0.addr == 8'h3E & write_0_en];	// <stdin>:3282:15, :3841:12, :3842:12, :3843:12, :3844:12, :3845:12, :3846:12, :3848:12
  assign _T_192 = Register_inst62;	// <stdin>:3848:12
  wire [31:0] _T_318 = ({{_T_191}, {write_0.data}})[write_0.addr == 8'h3F & write_0_en];	// <stdin>:3281:15, :3849:12, :3850:12, :3851:12, :3852:12, :3853:12, :3854:12, :3856:12
  assign _T_191 = Register_inst63;	// <stdin>:3856:12
  wire [31:0] _T_319 = ({{_T_190}, {write_0.data}})[write_0.addr == 8'h40 & write_0_en];	// <stdin>:3280:15, :3857:12, :3858:12, :3859:12, :3860:12, :3861:12, :3862:12, :3864:12
  assign _T_190 = Register_inst64;	// <stdin>:3864:12
  wire [31:0] _T_320 = ({{_T_189}, {write_0.data}})[write_0.addr == 8'h41 & write_0_en];	// <stdin>:3279:15, :3865:12, :3866:12, :3867:12, :3868:12, :3869:12, :3870:12, :3872:12
  assign _T_189 = Register_inst65;	// <stdin>:3872:12
  wire [31:0] _T_321 = ({{_T_188}, {write_0.data}})[write_0.addr == 8'h42 & write_0_en];	// <stdin>:3278:15, :3873:12, :3874:12, :3875:12, :3876:12, :3877:12, :3878:12, :3880:12
  assign _T_188 = Register_inst66;	// <stdin>:3880:12
  wire [31:0] _T_322 = ({{_T_187}, {write_0.data}})[write_0.addr == 8'h43 & write_0_en];	// <stdin>:3277:15, :3881:12, :3882:12, :3883:12, :3884:12, :3885:12, :3886:12, :3888:12
  assign _T_187 = Register_inst67;	// <stdin>:3888:12
  wire [31:0] _T_323 = ({{_T_186}, {write_0.data}})[write_0.addr == 8'h44 & write_0_en];	// <stdin>:3276:15, :3889:12, :3890:12, :3891:12, :3892:12, :3893:12, :3894:12, :3896:12
  assign _T_186 = Register_inst68;	// <stdin>:3896:12
  wire [31:0] _T_324 = ({{_T_185}, {write_0.data}})[write_0.addr == 8'h45 & write_0_en];	// <stdin>:3275:15, :3897:12, :3898:12, :3899:12, :3900:12, :3901:12, :3902:12, :3904:12
  assign _T_185 = Register_inst69;	// <stdin>:3904:12
  wire [31:0] _T_325 = ({{_T_184}, {write_0.data}})[write_0.addr == 8'h46 & write_0_en];	// <stdin>:3274:15, :3905:12, :3906:12, :3907:12, :3908:12, :3909:12, :3910:12, :3912:12
  assign _T_184 = Register_inst70;	// <stdin>:3912:12
  wire [31:0] _T_326 = ({{_T_183}, {write_0.data}})[write_0.addr == 8'h47 & write_0_en];	// <stdin>:3273:15, :3913:12, :3914:12, :3915:12, :3916:12, :3917:12, :3918:12, :3920:12
  assign _T_183 = Register_inst71;	// <stdin>:3920:12
  wire [31:0] _T_327 = ({{_T_182}, {write_0.data}})[write_0.addr == 8'h48 & write_0_en];	// <stdin>:3272:15, :3921:12, :3922:12, :3923:12, :3924:12, :3925:12, :3926:12, :3928:12
  assign _T_182 = Register_inst72;	// <stdin>:3928:12
  wire [31:0] _T_328 = ({{_T_181}, {write_0.data}})[write_0.addr == 8'h49 & write_0_en];	// <stdin>:3271:15, :3929:12, :3930:12, :3931:12, :3932:12, :3933:12, :3934:12, :3936:12
  assign _T_181 = Register_inst73;	// <stdin>:3936:12
  wire [31:0] _T_329 = ({{_T_180}, {write_0.data}})[write_0.addr == 8'h4A & write_0_en];	// <stdin>:3270:15, :3937:12, :3938:12, :3939:12, :3940:12, :3941:12, :3942:12, :3944:12
  assign _T_180 = Register_inst74;	// <stdin>:3944:12
  wire [31:0] _T_330 = ({{_T_179}, {write_0.data}})[write_0.addr == 8'h4B & write_0_en];	// <stdin>:3269:15, :3945:12, :3946:12, :3947:12, :3948:12, :3949:12, :3950:12, :3952:12
  assign _T_179 = Register_inst75;	// <stdin>:3952:12
  wire [31:0] _T_331 = ({{_T_178}, {write_0.data}})[write_0.addr == 8'h4C & write_0_en];	// <stdin>:3268:15, :3953:12, :3954:12, :3955:12, :3956:12, :3957:12, :3958:12, :3960:12
  assign _T_178 = Register_inst76;	// <stdin>:3960:12
  wire [31:0] _T_332 = ({{_T_177}, {write_0.data}})[write_0.addr == 8'h4D & write_0_en];	// <stdin>:3267:15, :3961:12, :3962:12, :3963:12, :3964:12, :3965:12, :3966:12, :3968:12
  assign _T_177 = Register_inst77;	// <stdin>:3968:12
  wire [31:0] _T_333 = ({{_T_176}, {write_0.data}})[write_0.addr == 8'h4E & write_0_en];	// <stdin>:3266:15, :3969:12, :3970:12, :3971:12, :3972:12, :3973:12, :3974:12, :3976:12
  assign _T_176 = Register_inst78;	// <stdin>:3976:12
  wire [31:0] _T_334 = ({{_T_175}, {write_0.data}})[write_0.addr == 8'h4F & write_0_en];	// <stdin>:3265:15, :3977:12, :3978:12, :3979:12, :3980:12, :3981:12, :3982:12, :3984:12
  assign _T_175 = Register_inst79;	// <stdin>:3984:12
  wire [31:0] _T_335 = ({{_T_174}, {write_0.data}})[write_0.addr == 8'h50 & write_0_en];	// <stdin>:3264:15, :3985:12, :3986:12, :3987:12, :3988:12, :3989:12, :3990:12, :3992:12
  assign _T_174 = Register_inst80;	// <stdin>:3992:12
  wire [31:0] _T_336 = ({{_T_173}, {write_0.data}})[write_0.addr == 8'h51 & write_0_en];	// <stdin>:3263:15, :3993:12, :3994:12, :3995:12, :3996:12, :3997:12, :3998:12, :4000:12
  assign _T_173 = Register_inst81;	// <stdin>:4000:12
  wire [31:0] _T_337 = ({{_T_172}, {write_0.data}})[write_0.addr == 8'h52 & write_0_en];	// <stdin>:3262:15, :4001:12, :4002:12, :4003:12, :4004:12, :4005:12, :4006:12, :4008:12
  assign _T_172 = Register_inst82;	// <stdin>:4008:12
  wire [31:0] _T_338 = ({{_T_171}, {write_0.data}})[write_0.addr == 8'h53 & write_0_en];	// <stdin>:3261:15, :4009:12, :4010:12, :4011:12, :4012:12, :4013:12, :4014:12, :4016:12
  assign _T_171 = Register_inst83;	// <stdin>:4016:12
  wire [31:0] _T_339 = ({{_T_170}, {write_0.data}})[write_0.addr == 8'h54 & write_0_en];	// <stdin>:3260:15, :4017:12, :4018:12, :4019:12, :4020:12, :4021:12, :4022:12, :4024:12
  assign _T_170 = Register_inst84;	// <stdin>:4024:12
  wire [31:0] _T_340 = ({{_T_169}, {write_0.data}})[write_0.addr == 8'h55 & write_0_en];	// <stdin>:3259:15, :4025:12, :4026:12, :4027:12, :4028:12, :4029:12, :4030:12, :4032:12
  assign _T_169 = Register_inst85;	// <stdin>:4032:12
  wire [31:0] _T_341 = ({{_T_168}, {write_0.data}})[write_0.addr == 8'h56 & write_0_en];	// <stdin>:3258:15, :4033:12, :4034:12, :4035:12, :4036:12, :4037:12, :4038:12, :4040:12
  assign _T_168 = Register_inst86;	// <stdin>:4040:12
  wire [31:0] _T_342 = ({{_T_167}, {write_0.data}})[write_0.addr == 8'h57 & write_0_en];	// <stdin>:3257:15, :4041:12, :4042:12, :4043:12, :4044:12, :4045:12, :4046:12, :4048:12
  assign _T_167 = Register_inst87;	// <stdin>:4048:12
  wire [31:0] _T_343 = ({{_T_166}, {write_0.data}})[write_0.addr == 8'h58 & write_0_en];	// <stdin>:3256:15, :4049:12, :4050:12, :4051:12, :4052:12, :4053:12, :4054:12, :4056:12
  assign _T_166 = Register_inst88;	// <stdin>:4056:12
  wire [31:0] _T_344 = ({{_T_165}, {write_0.data}})[write_0.addr == 8'h59 & write_0_en];	// <stdin>:3255:15, :4057:12, :4058:12, :4059:12, :4060:12, :4061:12, :4062:12, :4064:12
  assign _T_165 = Register_inst89;	// <stdin>:4064:12
  wire [31:0] _T_345 = ({{_T_164}, {write_0.data}})[write_0.addr == 8'h5A & write_0_en];	// <stdin>:3254:15, :4065:12, :4066:12, :4067:12, :4068:12, :4069:12, :4070:12, :4072:12
  assign _T_164 = Register_inst90;	// <stdin>:4072:12
  wire [31:0] _T_346 = ({{_T_163}, {write_0.data}})[write_0.addr == 8'h5B & write_0_en];	// <stdin>:3253:15, :4073:12, :4074:12, :4075:12, :4076:12, :4077:12, :4078:12, :4080:12
  assign _T_163 = Register_inst91;	// <stdin>:4080:12
  wire [31:0] _T_347 = ({{_T_162}, {write_0.data}})[write_0.addr == 8'h5C & write_0_en];	// <stdin>:3252:15, :4081:12, :4082:12, :4083:12, :4084:12, :4085:12, :4086:12, :4088:12
  assign _T_162 = Register_inst92;	// <stdin>:4088:12
  wire [31:0] _T_348 = ({{_T_161}, {write_0.data}})[write_0.addr == 8'h5D & write_0_en];	// <stdin>:3251:15, :4089:12, :4090:12, :4091:12, :4092:12, :4093:12, :4094:12, :4096:12
  assign _T_161 = Register_inst93;	// <stdin>:4096:12
  wire [31:0] _T_349 = ({{_T_160}, {write_0.data}})[write_0.addr == 8'h5E & write_0_en];	// <stdin>:3250:15, :4097:12, :4098:12, :4099:12, :4100:12, :4101:12, :4102:12, :4104:12
  assign _T_160 = Register_inst94;	// <stdin>:4104:12
  wire [31:0] _T_350 = ({{_T_159}, {write_0.data}})[write_0.addr == 8'h5F & write_0_en];	// <stdin>:3249:15, :4105:12, :4106:12, :4107:12, :4108:12, :4109:12, :4110:12, :4112:12
  assign _T_159 = Register_inst95;	// <stdin>:4112:12
  wire [31:0] _T_351 = ({{_T_158}, {write_0.data}})[write_0.addr == 8'h60 & write_0_en];	// <stdin>:3248:15, :4113:12, :4114:12, :4115:12, :4116:12, :4117:12, :4118:12, :4120:12
  assign _T_158 = Register_inst96;	// <stdin>:4120:12
  wire [31:0] _T_352 = ({{_T_157}, {write_0.data}})[write_0.addr == 8'h61 & write_0_en];	// <stdin>:3247:15, :4121:12, :4122:12, :4123:12, :4124:12, :4125:12, :4126:12, :4128:12
  assign _T_157 = Register_inst97;	// <stdin>:4128:12
  wire [31:0] _T_353 = ({{_T_156}, {write_0.data}})[write_0.addr == 8'h62 & write_0_en];	// <stdin>:3246:15, :4129:12, :4130:12, :4131:12, :4132:12, :4133:12, :4134:12, :4136:12
  assign _T_156 = Register_inst98;	// <stdin>:4136:12
  wire [31:0] _T_354 = ({{_T_155}, {write_0.data}})[write_0.addr == 8'h63 & write_0_en];	// <stdin>:3245:15, :4137:12, :4138:12, :4139:12, :4140:12, :4141:12, :4142:12, :4144:12
  assign _T_155 = Register_inst99;	// <stdin>:4144:12
  wire [31:0] _T_355 = ({{_T_154}, {write_0.data}})[write_0.addr == 8'h64 & write_0_en];	// <stdin>:3244:16, :4145:12, :4146:12, :4147:12, :4148:12, :4149:12, :4150:12, :4152:12
  assign _T_154 = Register_inst100;	// <stdin>:4152:12
  wire [31:0] _T_356 = ({{_T_153}, {write_0.data}})[write_0.addr == 8'h65 & write_0_en];	// <stdin>:3243:16, :4153:12, :4154:12, :4155:12, :4156:12, :4157:12, :4158:12, :4160:12
  assign _T_153 = Register_inst101;	// <stdin>:4160:12
  wire [31:0] _T_357 = ({{_T_152}, {write_0.data}})[write_0.addr == 8'h66 & write_0_en];	// <stdin>:3242:16, :4161:12, :4162:12, :4163:12, :4164:12, :4165:12, :4166:12, :4168:12
  assign _T_152 = Register_inst102;	// <stdin>:4168:12
  wire [31:0] _T_358 = ({{_T_151}, {write_0.data}})[write_0.addr == 8'h67 & write_0_en];	// <stdin>:3241:16, :4169:12, :4170:12, :4171:12, :4172:12, :4173:12, :4174:12, :4176:12
  assign _T_151 = Register_inst103;	// <stdin>:4176:12
  wire [31:0] _T_359 = ({{_T_150}, {write_0.data}})[write_0.addr == 8'h68 & write_0_en];	// <stdin>:3240:16, :4177:12, :4178:12, :4179:12, :4180:12, :4181:12, :4182:12, :4184:12
  assign _T_150 = Register_inst104;	// <stdin>:4184:12
  wire [31:0] _T_360 = ({{_T_149}, {write_0.data}})[write_0.addr == 8'h69 & write_0_en];	// <stdin>:3239:16, :4185:12, :4186:12, :4187:12, :4188:12, :4189:12, :4190:12, :4192:12
  assign _T_149 = Register_inst105;	// <stdin>:4192:12
  wire [31:0] _T_361 = ({{_T_148}, {write_0.data}})[write_0.addr == 8'h6A & write_0_en];	// <stdin>:3238:16, :4193:12, :4194:12, :4195:12, :4196:12, :4197:12, :4198:12, :4200:12
  assign _T_148 = Register_inst106;	// <stdin>:4200:12
  wire [31:0] _T_362 = ({{_T_147}, {write_0.data}})[write_0.addr == 8'h6B & write_0_en];	// <stdin>:3237:16, :4201:12, :4202:12, :4203:12, :4204:12, :4205:12, :4206:12, :4208:12
  assign _T_147 = Register_inst107;	// <stdin>:4208:12
  wire [31:0] _T_363 = ({{_T_146}, {write_0.data}})[write_0.addr == 8'h6C & write_0_en];	// <stdin>:3236:16, :4209:12, :4210:12, :4211:12, :4212:12, :4213:12, :4214:12, :4216:12
  assign _T_146 = Register_inst108;	// <stdin>:4216:12
  wire [31:0] _T_364 = ({{_T_145}, {write_0.data}})[write_0.addr == 8'h6D & write_0_en];	// <stdin>:3235:16, :4217:12, :4218:12, :4219:12, :4220:12, :4221:12, :4222:12, :4224:12
  assign _T_145 = Register_inst109;	// <stdin>:4224:12
  wire [31:0] _T_365 = ({{_T_144}, {write_0.data}})[write_0.addr == 8'h6E & write_0_en];	// <stdin>:3234:16, :4225:12, :4226:12, :4227:12, :4228:12, :4229:12, :4230:12, :4232:12
  assign _T_144 = Register_inst110;	// <stdin>:4232:12
  wire [31:0] _T_366 = ({{_T_143}, {write_0.data}})[write_0.addr == 8'h6F & write_0_en];	// <stdin>:3233:16, :4233:12, :4234:12, :4235:12, :4236:12, :4237:12, :4238:12, :4240:12
  assign _T_143 = Register_inst111;	// <stdin>:4240:12
  wire [31:0] _T_367 = ({{_T_142}, {write_0.data}})[write_0.addr == 8'h70 & write_0_en];	// <stdin>:3232:16, :4241:12, :4242:12, :4243:12, :4244:12, :4245:12, :4246:12, :4248:12
  assign _T_142 = Register_inst112;	// <stdin>:4248:12
  wire [31:0] _T_368 = ({{_T_141}, {write_0.data}})[write_0.addr == 8'h71 & write_0_en];	// <stdin>:3231:16, :4249:12, :4250:12, :4251:12, :4252:12, :4253:12, :4254:12, :4256:12
  assign _T_141 = Register_inst113;	// <stdin>:4256:12
  wire [31:0] _T_369 = ({{_T_140}, {write_0.data}})[write_0.addr == 8'h72 & write_0_en];	// <stdin>:3230:16, :4257:12, :4258:12, :4259:12, :4260:12, :4261:12, :4262:12, :4264:12
  assign _T_140 = Register_inst114;	// <stdin>:4264:12
  wire [31:0] _T_370 = ({{_T_139}, {write_0.data}})[write_0.addr == 8'h73 & write_0_en];	// <stdin>:3229:16, :4265:12, :4266:12, :4267:12, :4268:12, :4269:12, :4270:12, :4272:12
  assign _T_139 = Register_inst115;	// <stdin>:4272:12
  wire [31:0] _T_371 = ({{_T_138}, {write_0.data}})[write_0.addr == 8'h74 & write_0_en];	// <stdin>:3228:16, :4273:12, :4274:12, :4275:12, :4276:12, :4277:12, :4278:12, :4280:12
  assign _T_138 = Register_inst116;	// <stdin>:4280:12
  wire [31:0] _T_372 = ({{_T_137}, {write_0.data}})[write_0.addr == 8'h75 & write_0_en];	// <stdin>:3227:16, :4281:12, :4282:12, :4283:12, :4284:12, :4285:12, :4286:12, :4288:12
  assign _T_137 = Register_inst117;	// <stdin>:4288:12
  wire [31:0] _T_373 = ({{_T_136}, {write_0.data}})[write_0.addr == 8'h76 & write_0_en];	// <stdin>:3226:16, :4289:12, :4290:12, :4291:12, :4292:12, :4293:12, :4294:12, :4296:12
  assign _T_136 = Register_inst118;	// <stdin>:4296:12
  wire [31:0] _T_374 = ({{_T_135}, {write_0.data}})[write_0.addr == 8'h77 & write_0_en];	// <stdin>:3225:16, :4297:12, :4298:12, :4299:12, :4300:12, :4301:12, :4302:12, :4304:12
  assign _T_135 = Register_inst119;	// <stdin>:4304:12
  wire [31:0] _T_375 = ({{_T_134}, {write_0.data}})[write_0.addr == 8'h78 & write_0_en];	// <stdin>:3224:16, :4305:12, :4306:12, :4307:12, :4308:12, :4309:12, :4310:12, :4312:12
  assign _T_134 = Register_inst120;	// <stdin>:4312:12
  wire [31:0] _T_376 = ({{_T_133}, {write_0.data}})[write_0.addr == 8'h79 & write_0_en];	// <stdin>:3223:16, :4313:12, :4314:12, :4315:12, :4316:12, :4317:12, :4318:12, :4320:12
  assign _T_133 = Register_inst121;	// <stdin>:4320:12
  wire [31:0] _T_377 = ({{_T_132}, {write_0.data}})[write_0.addr == 8'h7A & write_0_en];	// <stdin>:3222:16, :4321:12, :4322:12, :4323:12, :4324:12, :4325:12, :4326:12, :4328:12
  assign _T_132 = Register_inst122;	// <stdin>:4328:12
  wire [31:0] _T_378 = ({{_T_131}, {write_0.data}})[write_0.addr == 8'h7B & write_0_en];	// <stdin>:3221:16, :4329:12, :4330:12, :4331:12, :4332:12, :4333:12, :4334:12, :4336:12
  assign _T_131 = Register_inst123;	// <stdin>:4336:12
  wire [31:0] _T_379 = ({{_T_130}, {write_0.data}})[write_0.addr == 8'h7C & write_0_en];	// <stdin>:3220:16, :4337:12, :4338:12, :4339:12, :4340:12, :4341:12, :4342:12, :4344:12
  assign _T_130 = Register_inst124;	// <stdin>:4344:12
  wire [31:0] _T_380 = ({{_T_129}, {write_0.data}})[write_0.addr == 8'h7D & write_0_en];	// <stdin>:3219:16, :4345:12, :4346:12, :4347:12, :4348:12, :4349:12, :4350:12, :4352:12
  assign _T_129 = Register_inst125;	// <stdin>:4352:12
  wire [31:0] _T_381 = ({{_T_128}, {write_0.data}})[write_0.addr == 8'h7E & write_0_en];	// <stdin>:3218:16, :4353:12, :4354:12, :4355:12, :4356:12, :4357:12, :4358:12, :4360:12
  assign _T_128 = Register_inst126;	// <stdin>:4360:12
  wire [31:0] _T_382 = ({{_T_127}, {write_0.data}})[write_0.addr == 8'h7F & write_0_en];	// <stdin>:3217:16, :4361:12, :4362:12, :4363:12, :4364:12, :4365:12, :4366:12, :4368:12
  assign _T_127 = Register_inst127;	// <stdin>:4368:12
  wire [31:0] _T_383 = ({{_T_126}, {write_0.data}})[write_0.addr == 8'h80 & write_0_en];	// <stdin>:3216:17, :4369:12, :4370:12, :4371:12, :4372:12, :4373:12, :4374:12, :4376:12
  assign _T_126 = Register_inst128;	// <stdin>:4376:12
  wire [31:0] _T_384 = ({{_T_125}, {write_0.data}})[write_0.addr == 8'h81 & write_0_en];	// <stdin>:3215:17, :4377:12, :4378:12, :4379:12, :4380:12, :4381:12, :4382:12, :4384:12
  assign _T_125 = Register_inst129;	// <stdin>:4384:12
  wire [31:0] _T_385 = ({{_T_124}, {write_0.data}})[write_0.addr == 8'h82 & write_0_en];	// <stdin>:3214:17, :4385:12, :4386:12, :4387:12, :4388:12, :4389:12, :4390:12, :4392:12
  assign _T_124 = Register_inst130;	// <stdin>:4392:12
  wire [31:0] _T_386 = ({{_T_123}, {write_0.data}})[write_0.addr == 8'h83 & write_0_en];	// <stdin>:3213:17, :4393:12, :4394:12, :4395:12, :4396:12, :4397:12, :4398:12, :4400:12
  assign _T_123 = Register_inst131;	// <stdin>:4400:12
  wire [31:0] _T_387 = ({{_T_122}, {write_0.data}})[write_0.addr == 8'h84 & write_0_en];	// <stdin>:3212:17, :4401:12, :4402:12, :4403:12, :4404:12, :4405:12, :4406:12, :4408:12
  assign _T_122 = Register_inst132;	// <stdin>:4408:12
  wire [31:0] _T_388 = ({{_T_121}, {write_0.data}})[write_0.addr == 8'h85 & write_0_en];	// <stdin>:3211:17, :4409:12, :4410:12, :4411:12, :4412:12, :4413:12, :4414:12, :4416:12
  assign _T_121 = Register_inst133;	// <stdin>:4416:12
  wire [31:0] _T_389 = ({{_T_120}, {write_0.data}})[write_0.addr == 8'h86 & write_0_en];	// <stdin>:3210:17, :4417:12, :4418:12, :4419:12, :4420:12, :4421:12, :4422:12, :4424:12
  assign _T_120 = Register_inst134;	// <stdin>:4424:12
  wire [31:0] _T_390 = ({{_T_119}, {write_0.data}})[write_0.addr == 8'h87 & write_0_en];	// <stdin>:3209:17, :4425:12, :4426:12, :4427:12, :4428:12, :4429:12, :4430:12, :4432:12
  assign _T_119 = Register_inst135;	// <stdin>:4432:12
  wire [31:0] _T_391 = ({{_T_118}, {write_0.data}})[write_0.addr == 8'h88 & write_0_en];	// <stdin>:3208:17, :4433:12, :4434:12, :4435:12, :4436:12, :4437:12, :4438:12, :4440:12
  assign _T_118 = Register_inst136;	// <stdin>:4440:12
  wire [31:0] _T_392 = ({{_T_117}, {write_0.data}})[write_0.addr == 8'h89 & write_0_en];	// <stdin>:3207:17, :4441:12, :4442:12, :4443:12, :4444:12, :4445:12, :4446:12, :4448:12
  assign _T_117 = Register_inst137;	// <stdin>:4448:12
  wire [31:0] _T_393 = ({{_T_116}, {write_0.data}})[write_0.addr == 8'h8A & write_0_en];	// <stdin>:3206:17, :4449:12, :4450:12, :4451:12, :4452:12, :4453:12, :4454:12, :4456:12
  assign _T_116 = Register_inst138;	// <stdin>:4456:12
  wire [31:0] _T_394 = ({{_T_115}, {write_0.data}})[write_0.addr == 8'h8B & write_0_en];	// <stdin>:3205:17, :4457:12, :4458:12, :4459:12, :4460:12, :4461:12, :4462:12, :4464:12
  assign _T_115 = Register_inst139;	// <stdin>:4464:12
  wire [31:0] _T_395 = ({{_T_114}, {write_0.data}})[write_0.addr == 8'h8C & write_0_en];	// <stdin>:3204:17, :4465:12, :4466:12, :4467:12, :4468:12, :4469:12, :4470:12, :4472:12
  assign _T_114 = Register_inst140;	// <stdin>:4472:12
  wire [31:0] _T_396 = ({{_T_113}, {write_0.data}})[write_0.addr == 8'h8D & write_0_en];	// <stdin>:3203:17, :4473:12, :4474:12, :4475:12, :4476:12, :4477:12, :4478:12, :4480:12
  assign _T_113 = Register_inst141;	// <stdin>:4480:12
  wire [31:0] _T_397 = ({{_T_112}, {write_0.data}})[write_0.addr == 8'h8E & write_0_en];	// <stdin>:3202:17, :4481:12, :4482:12, :4483:12, :4484:12, :4485:12, :4486:12, :4488:13
  assign _T_112 = Register_inst142;	// <stdin>:4488:13
  wire [31:0] _T_398 = ({{_T_111}, {write_0.data}})[write_0.addr == 8'h8F & write_0_en];	// <stdin>:3201:17, :4489:13, :4490:13, :4491:13, :4492:13, :4493:13, :4494:13, :4496:13
  assign _T_111 = Register_inst143;	// <stdin>:4496:13
  wire [31:0] _T_399 = ({{_T_110}, {write_0.data}})[write_0.addr == 8'h90 & write_0_en];	// <stdin>:3200:17, :4497:13, :4498:13, :4499:13, :4500:13, :4501:13, :4502:13, :4504:13
  assign _T_110 = Register_inst144;	// <stdin>:4504:13
  wire [31:0] _T_400 = ({{_T_109}, {write_0.data}})[write_0.addr == 8'h91 & write_0_en];	// <stdin>:3199:17, :4505:13, :4506:13, :4507:13, :4508:13, :4509:13, :4510:13, :4512:13
  assign _T_109 = Register_inst145;	// <stdin>:4512:13
  wire [31:0] _T_401 = ({{_T_108}, {write_0.data}})[write_0.addr == 8'h92 & write_0_en];	// <stdin>:3198:17, :4513:13, :4514:13, :4515:13, :4516:13, :4517:13, :4518:13, :4520:13
  assign _T_108 = Register_inst146;	// <stdin>:4520:13
  wire [31:0] _T_402 = ({{_T_107}, {write_0.data}})[write_0.addr == 8'h93 & write_0_en];	// <stdin>:3197:17, :4521:13, :4522:13, :4523:13, :4524:13, :4525:13, :4526:13, :4528:13
  assign _T_107 = Register_inst147;	// <stdin>:4528:13
  wire [31:0] _T_403 = ({{_T_106}, {write_0.data}})[write_0.addr == 8'h94 & write_0_en];	// <stdin>:3196:17, :4529:13, :4530:13, :4531:13, :4532:13, :4533:13, :4534:13, :4536:13
  assign _T_106 = Register_inst148;	// <stdin>:4536:13
  wire [31:0] _T_404 = ({{_T_105}, {write_0.data}})[write_0.addr == 8'h95 & write_0_en];	// <stdin>:3195:17, :4537:13, :4538:13, :4539:13, :4540:13, :4541:13, :4542:13, :4544:13
  assign _T_105 = Register_inst149;	// <stdin>:4544:13
  wire [31:0] _T_405 = ({{_T_104}, {write_0.data}})[write_0.addr == 8'h96 & write_0_en];	// <stdin>:3194:17, :4545:13, :4546:13, :4547:13, :4548:13, :4549:13, :4550:13, :4552:13
  assign _T_104 = Register_inst150;	// <stdin>:4552:13
  wire [31:0] _T_406 = ({{_T_103}, {write_0.data}})[write_0.addr == 8'h97 & write_0_en];	// <stdin>:3193:17, :4553:13, :4554:13, :4555:13, :4556:13, :4557:13, :4558:13, :4560:13
  assign _T_103 = Register_inst151;	// <stdin>:4560:13
  wire [31:0] _T_407 = ({{_T_102}, {write_0.data}})[write_0.addr == 8'h98 & write_0_en];	// <stdin>:3192:17, :4561:13, :4562:13, :4563:13, :4564:13, :4565:13, :4566:13, :4568:13
  assign _T_102 = Register_inst152;	// <stdin>:4568:13
  wire [31:0] _T_408 = ({{_T_101}, {write_0.data}})[write_0.addr == 8'h99 & write_0_en];	// <stdin>:3191:17, :4569:13, :4570:13, :4571:13, :4572:13, :4573:13, :4574:13, :4576:13
  assign _T_101 = Register_inst153;	// <stdin>:4576:13
  wire [31:0] _T_409 = ({{_T_100}, {write_0.data}})[write_0.addr == 8'h9A & write_0_en];	// <stdin>:3190:17, :4577:13, :4578:13, :4579:13, :4580:13, :4581:13, :4582:13, :4584:13
  assign _T_100 = Register_inst154;	// <stdin>:4584:13
  wire [31:0] _T_410 = ({{_T_99}, {write_0.data}})[write_0.addr == 8'h9B & write_0_en];	// <stdin>:3189:17, :4585:13, :4586:13, :4587:13, :4588:13, :4589:13, :4590:13, :4592:13
  assign _T_99 = Register_inst155;	// <stdin>:4592:13
  wire [31:0] _T_411 = ({{_T_98}, {write_0.data}})[write_0.addr == 8'h9C & write_0_en];	// <stdin>:3188:17, :4593:13, :4594:13, :4595:13, :4596:13, :4597:13, :4598:13, :4600:13
  assign _T_98 = Register_inst156;	// <stdin>:4600:13
  wire [31:0] _T_412 = ({{_T_97}, {write_0.data}})[write_0.addr == 8'h9D & write_0_en];	// <stdin>:3187:16, :4601:13, :4602:13, :4603:13, :4604:13, :4605:13, :4606:13, :4608:13
  assign _T_97 = Register_inst157;	// <stdin>:4608:13
  wire [31:0] _T_413 = ({{_T_96}, {write_0.data}})[write_0.addr == 8'h9E & write_0_en];	// <stdin>:3186:16, :4609:13, :4610:13, :4611:13, :4612:13, :4613:13, :4614:13, :4616:13
  assign _T_96 = Register_inst158;	// <stdin>:4616:13
  wire [31:0] _T_414 = ({{_T_95}, {write_0.data}})[write_0.addr == 8'h9F & write_0_en];	// <stdin>:3185:16, :4617:13, :4618:13, :4619:13, :4620:13, :4621:13, :4622:13, :4624:13
  assign _T_95 = Register_inst159;	// <stdin>:4624:13
  wire [31:0] _T_415 = ({{_T_94}, {write_0.data}})[write_0.addr == 8'hA0 & write_0_en];	// <stdin>:3184:16, :4625:13, :4626:13, :4627:13, :4628:13, :4629:13, :4630:13, :4632:13
  assign _T_94 = Register_inst160;	// <stdin>:4632:13
  wire [31:0] _T_416 = ({{_T_93}, {write_0.data}})[write_0.addr == 8'hA1 & write_0_en];	// <stdin>:3183:16, :4633:13, :4634:13, :4635:13, :4636:13, :4637:13, :4638:13, :4640:13
  assign _T_93 = Register_inst161;	// <stdin>:4640:13
  wire [31:0] _T_417 = ({{_T_92}, {write_0.data}})[write_0.addr == 8'hA2 & write_0_en];	// <stdin>:3182:16, :4641:13, :4642:13, :4643:13, :4644:13, :4645:13, :4646:13, :4648:13
  assign _T_92 = Register_inst162;	// <stdin>:4648:13
  wire [31:0] _T_418 = ({{_T_91}, {write_0.data}})[write_0.addr == 8'hA3 & write_0_en];	// <stdin>:3181:16, :4649:13, :4650:13, :4651:13, :4652:13, :4653:13, :4654:13, :4656:13
  assign _T_91 = Register_inst163;	// <stdin>:4656:13
  wire [31:0] _T_419 = ({{_T_90}, {write_0.data}})[write_0.addr == 8'hA4 & write_0_en];	// <stdin>:3180:16, :4657:13, :4658:13, :4659:13, :4660:13, :4661:13, :4662:13, :4664:13
  assign _T_90 = Register_inst164;	// <stdin>:4664:13
  wire [31:0] _T_420 = ({{_T_89}, {write_0.data}})[write_0.addr == 8'hA5 & write_0_en];	// <stdin>:3179:16, :4665:13, :4666:13, :4667:13, :4668:13, :4669:13, :4670:13, :4672:13
  assign _T_89 = Register_inst165;	// <stdin>:4672:13
  wire [31:0] _T_421 = ({{_T_88}, {write_0.data}})[write_0.addr == 8'hA6 & write_0_en];	// <stdin>:3178:16, :4673:13, :4674:13, :4675:13, :4676:13, :4677:13, :4678:13, :4680:13
  assign _T_88 = Register_inst166;	// <stdin>:4680:13
  wire [31:0] _T_422 = ({{_T_87}, {write_0.data}})[write_0.addr == 8'hA7 & write_0_en];	// <stdin>:3177:16, :4681:13, :4682:13, :4683:13, :4684:13, :4685:13, :4686:13, :4688:13
  assign _T_87 = Register_inst167;	// <stdin>:4688:13
  wire [31:0] _T_423 = ({{_T_86}, {write_0.data}})[write_0.addr == 8'hA8 & write_0_en];	// <stdin>:3176:16, :4689:13, :4690:13, :4691:13, :4692:13, :4693:13, :4694:13, :4696:13
  assign _T_86 = Register_inst168;	// <stdin>:4696:13
  wire [31:0] _T_424 = ({{_T_85}, {write_0.data}})[write_0.addr == 8'hA9 & write_0_en];	// <stdin>:3175:16, :4697:13, :4698:13, :4699:13, :4700:13, :4701:13, :4702:13, :4704:13
  assign _T_85 = Register_inst169;	// <stdin>:4704:13
  wire [31:0] _T_425 = ({{_T_84}, {write_0.data}})[write_0.addr == 8'hAA & write_0_en];	// <stdin>:3174:16, :4705:13, :4706:13, :4707:13, :4708:13, :4709:13, :4710:13, :4712:13
  assign _T_84 = Register_inst170;	// <stdin>:4712:13
  wire [31:0] _T_426 = ({{_T_83}, {write_0.data}})[write_0.addr == 8'hAB & write_0_en];	// <stdin>:3173:16, :4713:13, :4714:13, :4715:13, :4716:13, :4717:13, :4718:13, :4720:13
  assign _T_83 = Register_inst171;	// <stdin>:4720:13
  wire [31:0] _T_427 = ({{_T_82}, {write_0.data}})[write_0.addr == 8'hAC & write_0_en];	// <stdin>:3172:16, :4721:13, :4722:13, :4723:13, :4724:13, :4725:13, :4726:13, :4728:13
  assign _T_82 = Register_inst172;	// <stdin>:4728:13
  wire [31:0] _T_428 = ({{_T_81}, {write_0.data}})[write_0.addr == 8'hAD & write_0_en];	// <stdin>:3171:16, :4729:13, :4730:13, :4731:13, :4732:13, :4733:13, :4734:13, :4736:13
  assign _T_81 = Register_inst173;	// <stdin>:4736:13
  wire [31:0] _T_429 = ({{_T_80}, {write_0.data}})[write_0.addr == 8'hAE & write_0_en];	// <stdin>:3170:16, :4737:13, :4738:13, :4739:13, :4740:13, :4741:13, :4742:13, :4744:13
  assign _T_80 = Register_inst174;	// <stdin>:4744:13
  wire [31:0] _T_430 = ({{_T_79}, {write_0.data}})[write_0.addr == 8'hAF & write_0_en];	// <stdin>:3169:16, :4745:13, :4746:13, :4747:13, :4748:13, :4749:13, :4750:13, :4752:13
  assign _T_79 = Register_inst175;	// <stdin>:4752:13
  wire [31:0] _T_431 = ({{_T_78}, {write_0.data}})[write_0.addr == 8'hB0 & write_0_en];	// <stdin>:3168:16, :4753:13, :4754:13, :4755:13, :4756:13, :4757:13, :4758:13, :4760:13
  assign _T_78 = Register_inst176;	// <stdin>:4760:13
  wire [31:0] _T_432 = ({{_T_77}, {write_0.data}})[write_0.addr == 8'hB1 & write_0_en];	// <stdin>:3167:16, :4761:13, :4762:13, :4763:13, :4764:13, :4765:13, :4766:13, :4768:13
  assign _T_77 = Register_inst177;	// <stdin>:4768:13
  wire [31:0] _T_433 = ({{_T_76}, {write_0.data}})[write_0.addr == 8'hB2 & write_0_en];	// <stdin>:3166:16, :4769:13, :4770:13, :4771:13, :4772:13, :4773:13, :4774:13, :4776:13
  assign _T_76 = Register_inst178;	// <stdin>:4776:13
  wire [31:0] _T_434 = ({{_T_75}, {write_0.data}})[write_0.addr == 8'hB3 & write_0_en];	// <stdin>:3165:16, :4777:13, :4778:13, :4779:13, :4780:13, :4781:13, :4782:13, :4784:13
  assign _T_75 = Register_inst179;	// <stdin>:4784:13
  wire [31:0] _T_435 = ({{_T_74}, {write_0.data}})[write_0.addr == 8'hB4 & write_0_en];	// <stdin>:3164:16, :4785:13, :4786:13, :4787:13, :4788:13, :4789:13, :4790:13, :4792:13
  assign _T_74 = Register_inst180;	// <stdin>:4792:13
  wire [31:0] _T_436 = ({{_T_73}, {write_0.data}})[write_0.addr == 8'hB5 & write_0_en];	// <stdin>:3163:16, :4793:13, :4794:13, :4795:13, :4796:13, :4797:13, :4798:13, :4800:13
  assign _T_73 = Register_inst181;	// <stdin>:4800:13
  wire [31:0] _T_437 = ({{_T_72}, {write_0.data}})[write_0.addr == 8'hB6 & write_0_en];	// <stdin>:3162:16, :4801:13, :4802:13, :4803:13, :4804:13, :4805:13, :4806:13, :4808:13
  assign _T_72 = Register_inst182;	// <stdin>:4808:13
  wire [31:0] _T_438 = ({{_T_71}, {write_0.data}})[write_0.addr == 8'hB7 & write_0_en];	// <stdin>:3161:16, :4809:13, :4810:13, :4811:13, :4812:13, :4813:13, :4814:13, :4816:13
  assign _T_71 = Register_inst183;	// <stdin>:4816:13
  wire [31:0] _T_439 = ({{_T_70}, {write_0.data}})[write_0.addr == 8'hB8 & write_0_en];	// <stdin>:3160:16, :4817:13, :4818:13, :4819:13, :4820:13, :4821:13, :4822:13, :4824:13
  assign _T_70 = Register_inst184;	// <stdin>:4824:13
  wire [31:0] _T_440 = ({{_T_69}, {write_0.data}})[write_0.addr == 8'hB9 & write_0_en];	// <stdin>:3159:16, :4825:13, :4826:13, :4827:13, :4828:13, :4829:13, :4830:13, :4832:13
  assign _T_69 = Register_inst185;	// <stdin>:4832:13
  wire [31:0] _T_441 = ({{_T_68}, {write_0.data}})[write_0.addr == 8'hBA & write_0_en];	// <stdin>:3158:16, :4833:13, :4834:13, :4835:13, :4836:13, :4837:13, :4838:13, :4840:13
  assign _T_68 = Register_inst186;	// <stdin>:4840:13
  wire [31:0] _T_442 = ({{_T_67}, {write_0.data}})[write_0.addr == 8'hBB & write_0_en];	// <stdin>:3157:16, :4841:13, :4842:13, :4843:13, :4844:13, :4845:13, :4846:13, :4848:13
  assign _T_67 = Register_inst187;	// <stdin>:4848:13
  wire [31:0] _T_443 = ({{_T_66}, {write_0.data}})[write_0.addr == 8'hBC & write_0_en];	// <stdin>:3156:16, :4849:13, :4850:13, :4851:13, :4852:13, :4853:13, :4854:13, :4856:13
  assign _T_66 = Register_inst188;	// <stdin>:4856:13
  wire [31:0] _T_444 = ({{_T_65}, {write_0.data}})[write_0.addr == 8'hBD & write_0_en];	// <stdin>:3155:16, :4857:13, :4858:13, :4859:13, :4860:13, :4861:13, :4862:13, :4864:13
  assign _T_65 = Register_inst189;	// <stdin>:4864:13
  wire [31:0] _T_445 = ({{_T_64}, {write_0.data}})[write_0.addr == 8'hBE & write_0_en];	// <stdin>:3154:16, :4865:13, :4866:13, :4867:13, :4868:13, :4869:13, :4870:13, :4872:13
  assign _T_64 = Register_inst190;	// <stdin>:4872:13
  wire [31:0] _T_446 = ({{_T_63}, {write_0.data}})[write_0.addr == 8'hBF & write_0_en];	// <stdin>:3153:16, :4873:13, :4874:13, :4875:13, :4876:13, :4877:13, :4878:13, :4880:13
  assign _T_63 = Register_inst191;	// <stdin>:4880:13
  wire [31:0] _T_447 = ({{_T_62}, {write_0.data}})[write_0.addr == 8'hC0 & write_0_en];	// <stdin>:3152:16, :4881:13, :4882:13, :4883:13, :4884:13, :4885:13, :4886:13, :4888:13
  assign _T_62 = Register_inst192;	// <stdin>:4888:13
  wire [31:0] _T_448 = ({{_T_61}, {write_0.data}})[write_0.addr == 8'hC1 & write_0_en];	// <stdin>:3151:16, :4889:13, :4890:13, :4891:13, :4892:13, :4893:13, :4894:13, :4896:13
  assign _T_61 = Register_inst193;	// <stdin>:4896:13
  wire [31:0] _T_449 = ({{_T_60}, {write_0.data}})[write_0.addr == 8'hC2 & write_0_en];	// <stdin>:3150:16, :4897:13, :4898:13, :4899:13, :4900:13, :4901:13, :4902:13, :4904:13
  assign _T_60 = Register_inst194;	// <stdin>:4904:13
  wire [31:0] _T_450 = ({{_T_59}, {write_0.data}})[write_0.addr == 8'hC3 & write_0_en];	// <stdin>:3149:16, :4905:13, :4906:13, :4907:13, :4908:13, :4909:13, :4910:13, :4912:13
  assign _T_59 = Register_inst195;	// <stdin>:4912:13
  wire [31:0] _T_451 = ({{_T_58}, {write_0.data}})[write_0.addr == 8'hC4 & write_0_en];	// <stdin>:3148:16, :4913:13, :4914:13, :4915:13, :4916:13, :4917:13, :4918:13, :4920:13
  assign _T_58 = Register_inst196;	// <stdin>:4920:13
  wire [31:0] _T_452 = ({{_T_57}, {write_0.data}})[write_0.addr == 8'hC5 & write_0_en];	// <stdin>:3147:16, :4921:13, :4922:13, :4923:13, :4924:13, :4925:13, :4926:13, :4928:13
  assign _T_57 = Register_inst197;	// <stdin>:4928:13
  wire [31:0] _T_453 = ({{_T_56}, {write_0.data}})[write_0.addr == 8'hC6 & write_0_en];	// <stdin>:3146:16, :4929:13, :4930:13, :4931:13, :4932:13, :4933:13, :4934:13, :4936:13
  assign _T_56 = Register_inst198;	// <stdin>:4936:13
  wire [31:0] _T_454 = ({{_T_55}, {write_0.data}})[write_0.addr == 8'hC7 & write_0_en];	// <stdin>:3145:16, :4937:13, :4938:13, :4939:13, :4940:13, :4941:13, :4942:13, :4944:13
  assign _T_55 = Register_inst199;	// <stdin>:4944:13
  wire [31:0] _T_455 = ({{_T_54}, {write_0.data}})[write_0.addr == 8'hC8 & write_0_en];	// <stdin>:3144:16, :4945:13, :4946:13, :4947:13, :4948:13, :4949:13, :4950:13, :4952:13
  assign _T_54 = Register_inst200;	// <stdin>:4952:13
  wire [31:0] _T_456 = ({{_T_53}, {write_0.data}})[write_0.addr == 8'hC9 & write_0_en];	// <stdin>:3143:16, :4953:13, :4954:13, :4955:13, :4956:13, :4957:13, :4958:13, :4960:13
  assign _T_53 = Register_inst201;	// <stdin>:4960:13
  wire [31:0] _T_457 = ({{_T_52}, {write_0.data}})[write_0.addr == 8'hCA & write_0_en];	// <stdin>:3142:16, :4961:13, :4962:13, :4963:13, :4964:13, :4965:13, :4966:13, :4968:13
  assign _T_52 = Register_inst202;	// <stdin>:4968:13
  wire [31:0] _T_458 = ({{_T_51}, {write_0.data}})[write_0.addr == 8'hCB & write_0_en];	// <stdin>:3141:16, :4969:13, :4970:13, :4971:13, :4972:13, :4973:13, :4974:13, :4976:13
  assign _T_51 = Register_inst203;	// <stdin>:4976:13
  wire [31:0] _T_459 = ({{_T_50}, {write_0.data}})[write_0.addr == 8'hCC & write_0_en];	// <stdin>:3140:16, :4977:13, :4978:13, :4979:13, :4980:13, :4981:13, :4982:13, :4984:13
  assign _T_50 = Register_inst204;	// <stdin>:4984:13
  wire [31:0] _T_460 = ({{_T_49}, {write_0.data}})[write_0.addr == 8'hCD & write_0_en];	// <stdin>:3139:16, :4985:13, :4986:13, :4987:13, :4988:13, :4989:13, :4990:13, :4992:13
  assign _T_49 = Register_inst205;	// <stdin>:4992:13
  wire [31:0] _T_461 = ({{_T_48}, {write_0.data}})[write_0.addr == 8'hCE & write_0_en];	// <stdin>:3138:16, :4993:13, :4994:13, :4995:13, :4996:13, :4997:13, :4998:13, :5000:13
  assign _T_48 = Register_inst206;	// <stdin>:5000:13
  wire [31:0] _T_462 = ({{_T_47}, {write_0.data}})[write_0.addr == 8'hCF & write_0_en];	// <stdin>:3137:16, :5001:13, :5002:13, :5003:13, :5004:13, :5005:13, :5006:13, :5008:13
  assign _T_47 = Register_inst207;	// <stdin>:5008:13
  wire [31:0] _T_463 = ({{_T_46}, {write_0.data}})[write_0.addr == 8'hD0 & write_0_en];	// <stdin>:3136:16, :5009:13, :5010:13, :5011:13, :5012:13, :5013:13, :5014:13, :5016:13
  assign _T_46 = Register_inst208;	// <stdin>:5016:13
  wire [31:0] _T_464 = ({{_T_45}, {write_0.data}})[write_0.addr == 8'hD1 & write_0_en];	// <stdin>:3135:16, :5017:13, :5018:13, :5019:13, :5020:13, :5021:13, :5022:13, :5024:13
  assign _T_45 = Register_inst209;	// <stdin>:5024:13
  wire [31:0] _T_465 = ({{_T_44}, {write_0.data}})[write_0.addr == 8'hD2 & write_0_en];	// <stdin>:3134:16, :5025:13, :5026:13, :5027:13, :5028:13, :5029:13, :5030:13, :5032:13
  assign _T_44 = Register_inst210;	// <stdin>:5032:13
  wire [31:0] _T_466 = ({{_T_43}, {write_0.data}})[write_0.addr == 8'hD3 & write_0_en];	// <stdin>:3133:16, :5033:13, :5034:13, :5035:13, :5036:13, :5037:13, :5038:13, :5040:13
  assign _T_43 = Register_inst211;	// <stdin>:5040:13
  wire [31:0] _T_467 = ({{_T_42}, {write_0.data}})[write_0.addr == 8'hD4 & write_0_en];	// <stdin>:3132:16, :5041:13, :5042:13, :5043:13, :5044:13, :5045:13, :5046:13, :5048:13
  assign _T_42 = Register_inst212;	// <stdin>:5048:13
  wire [31:0] _T_468 = ({{_T_41}, {write_0.data}})[write_0.addr == 8'hD5 & write_0_en];	// <stdin>:3131:16, :5049:13, :5050:13, :5051:13, :5052:13, :5053:13, :5054:13, :5056:13
  assign _T_41 = Register_inst213;	// <stdin>:5056:13
  wire [31:0] _T_469 = ({{_T_40}, {write_0.data}})[write_0.addr == 8'hD6 & write_0_en];	// <stdin>:3130:16, :5057:13, :5058:13, :5059:13, :5060:13, :5061:13, :5062:13, :5064:13
  assign _T_40 = Register_inst214;	// <stdin>:5064:13
  wire [31:0] _T_470 = ({{_T_39}, {write_0.data}})[write_0.addr == 8'hD7 & write_0_en];	// <stdin>:3129:16, :5065:13, :5066:13, :5067:13, :5068:13, :5069:13, :5070:13, :5072:13
  assign _T_39 = Register_inst215;	// <stdin>:5072:13
  wire [31:0] _T_471 = ({{_T_38}, {write_0.data}})[write_0.addr == 8'hD8 & write_0_en];	// <stdin>:3128:16, :5073:13, :5074:13, :5075:13, :5076:13, :5077:13, :5078:13, :5080:13
  assign _T_38 = Register_inst216;	// <stdin>:5080:13
  wire [31:0] _T_472 = ({{_T_37}, {write_0.data}})[write_0.addr == 8'hD9 & write_0_en];	// <stdin>:3127:16, :5081:13, :5082:13, :5083:13, :5084:13, :5085:13, :5086:13, :5088:13
  assign _T_37 = Register_inst217;	// <stdin>:5088:13
  wire [31:0] _T_473 = ({{_T_36}, {write_0.data}})[write_0.addr == 8'hDA & write_0_en];	// <stdin>:3126:16, :5089:13, :5090:13, :5091:13, :5092:13, :5093:13, :5094:13, :5096:13
  assign _T_36 = Register_inst218;	// <stdin>:5096:13
  wire [31:0] _T_474 = ({{_T_35}, {write_0.data}})[write_0.addr == 8'hDB & write_0_en];	// <stdin>:3125:16, :5097:13, :5098:13, :5099:13, :5100:13, :5101:13, :5102:13, :5104:13
  assign _T_35 = Register_inst219;	// <stdin>:5104:13
  wire [31:0] _T_475 = ({{_T_34}, {write_0.data}})[write_0.addr == 8'hDC & write_0_en];	// <stdin>:3124:16, :5105:13, :5106:13, :5107:13, :5108:13, :5109:13, :5110:13, :5112:13
  assign _T_34 = Register_inst220;	// <stdin>:5112:13
  wire [31:0] _T_476 = ({{_T_33}, {write_0.data}})[write_0.addr == 8'hDD & write_0_en];	// <stdin>:3123:16, :5113:13, :5114:13, :5115:13, :5116:13, :5117:13, :5118:13, :5120:13
  assign _T_33 = Register_inst221;	// <stdin>:5120:13
  wire [31:0] _T_477 = ({{_T_32}, {write_0.data}})[write_0.addr == 8'hDE & write_0_en];	// <stdin>:3122:16, :5121:13, :5122:13, :5123:13, :5124:13, :5125:13, :5126:13, :5128:13
  assign _T_32 = Register_inst222;	// <stdin>:5128:13
  wire [31:0] _T_478 = ({{_T_31}, {write_0.data}})[write_0.addr == 8'hDF & write_0_en];	// <stdin>:3121:16, :5129:13, :5130:13, :5131:13, :5132:13, :5133:13, :5134:13, :5136:13
  assign _T_31 = Register_inst223;	// <stdin>:5136:13
  wire [31:0] _T_479 = ({{_T_30}, {write_0.data}})[write_0.addr == 8'hE0 & write_0_en];	// <stdin>:3120:16, :5137:13, :5138:13, :5139:13, :5140:13, :5141:13, :5142:13, :5144:13
  assign _T_30 = Register_inst224;	// <stdin>:5144:13
  wire [31:0] _T_480 = ({{_T_29}, {write_0.data}})[write_0.addr == 8'hE1 & write_0_en];	// <stdin>:3119:16, :5145:13, :5146:13, :5147:13, :5148:13, :5149:13, :5150:13, :5152:13
  assign _T_29 = Register_inst225;	// <stdin>:5152:13
  wire [31:0] _T_481 = ({{_T_28}, {write_0.data}})[write_0.addr == 8'hE2 & write_0_en];	// <stdin>:3118:16, :5153:13, :5154:13, :5155:13, :5156:13, :5157:13, :5158:13, :5160:13
  assign _T_28 = Register_inst226;	// <stdin>:5160:13
  wire [31:0] _T_482 = ({{_T_27}, {write_0.data}})[write_0.addr == 8'hE3 & write_0_en];	// <stdin>:3117:16, :5161:13, :5162:13, :5163:13, :5164:13, :5165:13, :5166:13, :5168:13
  assign _T_27 = Register_inst227;	// <stdin>:5168:13
  wire [31:0] _T_483 = ({{_T_26}, {write_0.data}})[write_0.addr == 8'hE4 & write_0_en];	// <stdin>:3116:16, :5169:13, :5170:13, :5171:13, :5172:13, :5173:13, :5174:13, :5176:13
  assign _T_26 = Register_inst228;	// <stdin>:5176:13
  wire [31:0] _T_484 = ({{_T_25}, {write_0.data}})[write_0.addr == 8'hE5 & write_0_en];	// <stdin>:3115:16, :5177:13, :5178:13, :5179:13, :5180:13, :5181:13, :5182:13, :5184:13
  assign _T_25 = Register_inst229;	// <stdin>:5184:13
  wire [31:0] _T_485 = ({{_T_24}, {write_0.data}})[write_0.addr == 8'hE6 & write_0_en];	// <stdin>:3114:16, :5185:13, :5186:13, :5187:13, :5188:13, :5189:13, :5190:13, :5192:13
  assign _T_24 = Register_inst230;	// <stdin>:5192:13
  wire [31:0] _T_486 = ({{_T_23}, {write_0.data}})[write_0.addr == 8'hE7 & write_0_en];	// <stdin>:3113:16, :5193:13, :5194:13, :5195:13, :5196:13, :5197:13, :5198:13, :5200:13
  assign _T_23 = Register_inst231;	// <stdin>:5200:13
  wire [31:0] _T_487 = ({{_T_22}, {write_0.data}})[write_0.addr == 8'hE8 & write_0_en];	// <stdin>:3112:16, :5201:13, :5202:13, :5203:13, :5204:13, :5205:13, :5206:13, :5208:13
  assign _T_22 = Register_inst232;	// <stdin>:5208:13
  wire [31:0] _T_488 = ({{_T_21}, {write_0.data}})[write_0.addr == 8'hE9 & write_0_en];	// <stdin>:3111:16, :5209:13, :5210:13, :5211:13, :5212:13, :5213:13, :5214:13, :5216:13
  assign _T_21 = Register_inst233;	// <stdin>:5216:13
  wire [31:0] _T_489 = ({{_T_20}, {write_0.data}})[write_0.addr == 8'hEA & write_0_en];	// <stdin>:3110:16, :5217:13, :5218:13, :5219:13, :5220:13, :5221:13, :5222:13, :5224:13
  assign _T_20 = Register_inst234;	// <stdin>:5224:13
  wire [31:0] _T_490 = ({{_T_19}, {write_0.data}})[write_0.addr == 8'hEB & write_0_en];	// <stdin>:3109:16, :5225:13, :5226:13, :5227:13, :5228:13, :5229:13, :5230:13, :5232:13
  assign _T_19 = Register_inst235;	// <stdin>:5232:13
  wire [31:0] _T_491 = ({{_T_18}, {write_0.data}})[write_0.addr == 8'hEC & write_0_en];	// <stdin>:3108:16, :5233:13, :5234:13, :5235:13, :5236:13, :5237:13, :5238:13, :5240:13
  assign _T_18 = Register_inst236;	// <stdin>:5240:13
  wire [31:0] _T_492 = ({{_T_17}, {write_0.data}})[write_0.addr == 8'hED & write_0_en];	// <stdin>:3107:16, :5241:13, :5242:13, :5243:13, :5244:13, :5245:13, :5246:13, :5248:13
  assign _T_17 = Register_inst237;	// <stdin>:5248:13
  wire [31:0] _T_493 = ({{_T_16}, {write_0.data}})[write_0.addr == 8'hEE & write_0_en];	// <stdin>:3106:16, :5249:13, :5250:13, :5251:13, :5252:13, :5253:13, :5254:13, :5256:13
  assign _T_16 = Register_inst238;	// <stdin>:5256:13
  wire [31:0] _T_494 = ({{_T_15}, {write_0.data}})[write_0.addr == 8'hEF & write_0_en];	// <stdin>:3105:16, :5257:13, :5258:13, :5259:13, :5260:13, :5261:13, :5262:13, :5264:13
  assign _T_15 = Register_inst239;	// <stdin>:5264:13
  wire [31:0] _T_495 = ({{_T_14}, {write_0.data}})[write_0.addr == 8'hF0 & write_0_en];	// <stdin>:3104:16, :5265:13, :5266:13, :5267:13, :5268:13, :5269:13, :5270:13, :5272:13
  assign _T_14 = Register_inst240;	// <stdin>:5272:13
  wire [31:0] _T_496 = ({{_T_13}, {write_0.data}})[write_0.addr == 8'hF1 & write_0_en];	// <stdin>:3103:16, :5273:13, :5274:13, :5275:13, :5276:13, :5277:13, :5278:13, :5280:13
  assign _T_13 = Register_inst241;	// <stdin>:5280:13
  wire [31:0] _T_497 = ({{_T_12}, {write_0.data}})[write_0.addr == 8'hF2 & write_0_en];	// <stdin>:3102:16, :5281:13, :5282:13, :5283:13, :5284:13, :5285:13, :5286:13, :5288:13
  assign _T_12 = Register_inst242;	// <stdin>:5288:13
  wire [31:0] _T_498 = ({{_T_11}, {write_0.data}})[write_0.addr == 8'hF3 & write_0_en];	// <stdin>:3101:16, :5289:13, :5290:13, :5291:13, :5292:13, :5293:13, :5294:13, :5296:13
  assign _T_11 = Register_inst243;	// <stdin>:5296:13
  wire [31:0] _T_499 = ({{_T_10}, {write_0.data}})[write_0.addr == 8'hF4 & write_0_en];	// <stdin>:3100:16, :5297:13, :5298:13, :5299:13, :5300:13, :5301:13, :5302:13, :5304:13
  assign _T_10 = Register_inst244;	// <stdin>:5304:13
  wire [31:0] _T_500 = ({{_T_9}, {write_0.data}})[write_0.addr == 8'hF5 & write_0_en];	// <stdin>:3099:16, :5305:13, :5306:13, :5307:13, :5308:13, :5309:13, :5310:13, :5312:13
  assign _T_9 = Register_inst245;	// <stdin>:5312:13
  wire [31:0] _T_501 = ({{_T_8}, {write_0.data}})[write_0.addr == 8'hF6 & write_0_en];	// <stdin>:3098:16, :5313:13, :5314:13, :5315:13, :5316:13, :5317:13, :5318:13, :5320:13
  assign _T_8 = Register_inst246;	// <stdin>:5320:13
  wire [31:0] _T_502 = ({{_T_7}, {write_0.data}})[write_0.addr == 8'hF7 & write_0_en];	// <stdin>:3097:15, :5321:13, :5322:13, :5323:13, :5324:13, :5325:13, :5326:13, :5328:13
  assign _T_7 = Register_inst247;	// <stdin>:5328:13
  wire [31:0] _T_503 = ({{_T_6}, {write_0.data}})[write_0.addr == 8'hF8 & write_0_en];	// <stdin>:3096:15, :5329:13, :5330:13, :5331:13, :5332:13, :5333:13, :5334:13, :5336:13
  assign _T_6 = Register_inst248;	// <stdin>:5336:13
  wire [31:0] _T_504 = ({{_T_5}, {write_0.data}})[write_0.addr == 8'hF9 & write_0_en];	// <stdin>:3095:15, :5337:13, :5338:13, :5339:13, :5340:13, :5341:13, :5342:13, :5344:13
  assign _T_5 = Register_inst249;	// <stdin>:5344:13
  wire [31:0] _T_505 = ({{_T_4}, {write_0.data}})[write_0.addr == 8'hFA & write_0_en];	// <stdin>:3094:15, :5345:13, :5346:13, :5347:13, :5348:13, :5349:13, :5350:13, :5352:13
  assign _T_4 = Register_inst250;	// <stdin>:5352:13
  wire [31:0] _T_506 = ({{_T_3}, {write_0.data}})[write_0.addr == 8'hFB & write_0_en];	// <stdin>:3093:15, :5353:13, :5354:13, :5355:13, :5356:13, :5357:13, :5358:13, :5360:13
  assign _T_3 = Register_inst251;	// <stdin>:5360:13
  wire [31:0] _T_507 = ({{_T_2}, {write_0.data}})[write_0.addr == 8'hFC & write_0_en];	// <stdin>:3092:15, :5361:13, :5362:13, :5363:13, :5364:13, :5365:13, :5366:13, :5368:13
  assign _T_2 = Register_inst252;	// <stdin>:5368:13
  wire [31:0] _T_508 = ({{_T_1}, {write_0.data}})[write_0.addr == 8'hFD & write_0_en];	// <stdin>:3091:15, :5369:13, :5370:13, :5371:13, :5372:13, :5373:13, :5374:13, :5376:13
  assign _T_1 = Register_inst253;	// <stdin>:5376:13
  wire [31:0] _T_509 = ({{_T_0}, {write_0.data}})[write_0.addr == 8'hFE & write_0_en];	// <stdin>:3090:15, :5377:13, :5378:13, :5379:13, :5380:13, :5381:13, :5382:13, :5384:13
  assign _T_0 = Register_inst254;	// <stdin>:5384:13
  wire [31:0] _T_510 = ({{_T}, {write_0.data}})[&write_0.addr & write_0_en];	// <stdin>:5385:13, :5386:13, :5387:13, :5388:13, :5389:13, :5390:13, :6167:13
  always @(posedge CLK or posedge ASYNCRESET) begin	// <stdin>:5392:5
    if (ASYNCRESET) begin	// <stdin>:5392:5
      Register_inst0 <= 32'h0;	// <stdin>:5650:17, :5651:7
      Register_inst1 <= 32'h0;	// <stdin>:5650:17, :5652:7
      Register_inst2 <= 32'h0;	// <stdin>:5650:17, :5653:7
      Register_inst3 <= 32'h0;	// <stdin>:5650:17, :5654:7
      Register_inst4 <= 32'h0;	// <stdin>:5650:17, :5655:7
      Register_inst5 <= 32'h0;	// <stdin>:5650:17, :5656:7
      Register_inst6 <= 32'h0;	// <stdin>:5650:17, :5657:7
      Register_inst7 <= 32'h0;	// <stdin>:5650:17, :5658:7
      Register_inst8 <= 32'h0;	// <stdin>:5650:17, :5659:7
      Register_inst9 <= 32'h0;	// <stdin>:5650:17, :5660:7
      Register_inst10 <= 32'h0;	// <stdin>:5650:17, :5661:7
      Register_inst11 <= 32'h0;	// <stdin>:5650:17, :5662:7
      Register_inst12 <= 32'h0;	// <stdin>:5650:17, :5663:7
      Register_inst13 <= 32'h0;	// <stdin>:5650:17, :5664:7
      Register_inst14 <= 32'h0;	// <stdin>:5650:17, :5665:7
      Register_inst15 <= 32'h0;	// <stdin>:5650:17, :5666:7
      Register_inst16 <= 32'h0;	// <stdin>:5650:17, :5667:7
      Register_inst17 <= 32'h0;	// <stdin>:5650:17, :5668:7
      Register_inst18 <= 32'h0;	// <stdin>:5650:17, :5669:7
      Register_inst19 <= 32'h0;	// <stdin>:5650:17, :5670:7
      Register_inst20 <= 32'h0;	// <stdin>:5650:17, :5671:7
      Register_inst21 <= 32'h0;	// <stdin>:5650:17, :5672:7
      Register_inst22 <= 32'h0;	// <stdin>:5650:17, :5673:7
      Register_inst23 <= 32'h0;	// <stdin>:5650:17, :5674:7
      Register_inst24 <= 32'h0;	// <stdin>:5650:17, :5675:7
      Register_inst25 <= 32'h0;	// <stdin>:5650:17, :5676:7
      Register_inst26 <= 32'h0;	// <stdin>:5650:17, :5677:7
      Register_inst27 <= 32'h0;	// <stdin>:5650:17, :5678:7
      Register_inst28 <= 32'h0;	// <stdin>:5650:17, :5679:7
      Register_inst29 <= 32'h0;	// <stdin>:5650:17, :5680:7
      Register_inst30 <= 32'h0;	// <stdin>:5650:17, :5681:7
      Register_inst31 <= 32'h0;	// <stdin>:5650:17, :5682:7
      Register_inst32 <= 32'h0;	// <stdin>:5650:17, :5683:7
      Register_inst33 <= 32'h0;	// <stdin>:5650:17, :5684:7
      Register_inst34 <= 32'h0;	// <stdin>:5650:17, :5685:7
      Register_inst35 <= 32'h0;	// <stdin>:5650:17, :5686:7
      Register_inst36 <= 32'h0;	// <stdin>:5650:17, :5687:7
      Register_inst37 <= 32'h0;	// <stdin>:5650:17, :5688:7
      Register_inst38 <= 32'h0;	// <stdin>:5650:17, :5689:7
      Register_inst39 <= 32'h0;	// <stdin>:5650:17, :5690:7
      Register_inst40 <= 32'h0;	// <stdin>:5650:17, :5691:7
      Register_inst41 <= 32'h0;	// <stdin>:5650:17, :5692:7
      Register_inst42 <= 32'h0;	// <stdin>:5650:17, :5693:7
      Register_inst43 <= 32'h0;	// <stdin>:5650:17, :5694:7
      Register_inst44 <= 32'h0;	// <stdin>:5650:17, :5695:7
      Register_inst45 <= 32'h0;	// <stdin>:5650:17, :5696:7
      Register_inst46 <= 32'h0;	// <stdin>:5650:17, :5697:7
      Register_inst47 <= 32'h0;	// <stdin>:5650:17, :5698:7
      Register_inst48 <= 32'h0;	// <stdin>:5650:17, :5699:7
      Register_inst49 <= 32'h0;	// <stdin>:5650:17, :5700:7
      Register_inst50 <= 32'h0;	// <stdin>:5650:17, :5701:7
      Register_inst51 <= 32'h0;	// <stdin>:5650:17, :5702:7
      Register_inst52 <= 32'h0;	// <stdin>:5650:17, :5703:7
      Register_inst53 <= 32'h0;	// <stdin>:5650:17, :5704:7
      Register_inst54 <= 32'h0;	// <stdin>:5650:17, :5705:7
      Register_inst55 <= 32'h0;	// <stdin>:5650:17, :5706:7
      Register_inst56 <= 32'h0;	// <stdin>:5650:17, :5707:7
      Register_inst57 <= 32'h0;	// <stdin>:5650:17, :5708:7
      Register_inst58 <= 32'h0;	// <stdin>:5650:17, :5709:7
      Register_inst59 <= 32'h0;	// <stdin>:5650:17, :5710:7
      Register_inst60 <= 32'h0;	// <stdin>:5650:17, :5711:7
      Register_inst61 <= 32'h0;	// <stdin>:5650:17, :5712:7
      Register_inst62 <= 32'h0;	// <stdin>:5650:17, :5713:7
      Register_inst63 <= 32'h0;	// <stdin>:5650:17, :5714:7
      Register_inst64 <= 32'h0;	// <stdin>:5650:17, :5715:7
      Register_inst65 <= 32'h0;	// <stdin>:5650:17, :5716:7
      Register_inst66 <= 32'h0;	// <stdin>:5650:17, :5717:7
      Register_inst67 <= 32'h0;	// <stdin>:5650:17, :5718:7
      Register_inst68 <= 32'h0;	// <stdin>:5650:17, :5719:7
      Register_inst69 <= 32'h0;	// <stdin>:5650:17, :5720:7
      Register_inst70 <= 32'h0;	// <stdin>:5650:17, :5721:7
      Register_inst71 <= 32'h0;	// <stdin>:5650:17, :5722:7
      Register_inst72 <= 32'h0;	// <stdin>:5650:17, :5723:7
      Register_inst73 <= 32'h0;	// <stdin>:5650:17, :5724:7
      Register_inst74 <= 32'h0;	// <stdin>:5650:17, :5725:7
      Register_inst75 <= 32'h0;	// <stdin>:5650:17, :5726:7
      Register_inst76 <= 32'h0;	// <stdin>:5650:17, :5727:7
      Register_inst77 <= 32'h0;	// <stdin>:5650:17, :5728:7
      Register_inst78 <= 32'h0;	// <stdin>:5650:17, :5729:7
      Register_inst79 <= 32'h0;	// <stdin>:5650:17, :5730:7
      Register_inst80 <= 32'h0;	// <stdin>:5650:17, :5731:7
      Register_inst81 <= 32'h0;	// <stdin>:5650:17, :5732:7
      Register_inst82 <= 32'h0;	// <stdin>:5650:17, :5733:7
      Register_inst83 <= 32'h0;	// <stdin>:5650:17, :5734:7
      Register_inst84 <= 32'h0;	// <stdin>:5650:17, :5735:7
      Register_inst85 <= 32'h0;	// <stdin>:5650:17, :5736:7
      Register_inst86 <= 32'h0;	// <stdin>:5650:17, :5737:7
      Register_inst87 <= 32'h0;	// <stdin>:5650:17, :5738:7
      Register_inst88 <= 32'h0;	// <stdin>:5650:17, :5739:7
      Register_inst89 <= 32'h0;	// <stdin>:5650:17, :5740:7
      Register_inst90 <= 32'h0;	// <stdin>:5650:17, :5741:7
      Register_inst91 <= 32'h0;	// <stdin>:5650:17, :5742:7
      Register_inst92 <= 32'h0;	// <stdin>:5650:17, :5743:7
      Register_inst93 <= 32'h0;	// <stdin>:5650:17, :5744:7
      Register_inst94 <= 32'h0;	// <stdin>:5650:17, :5745:7
      Register_inst95 <= 32'h0;	// <stdin>:5650:17, :5746:7
      Register_inst96 <= 32'h0;	// <stdin>:5650:17, :5747:7
      Register_inst97 <= 32'h0;	// <stdin>:5650:17, :5748:7
      Register_inst98 <= 32'h0;	// <stdin>:5650:17, :5749:7
      Register_inst99 <= 32'h0;	// <stdin>:5650:17, :5750:7
      Register_inst100 <= 32'h0;	// <stdin>:5650:17, :5751:7
      Register_inst101 <= 32'h0;	// <stdin>:5650:17, :5752:7
      Register_inst102 <= 32'h0;	// <stdin>:5650:17, :5753:7
      Register_inst103 <= 32'h0;	// <stdin>:5650:17, :5754:7
      Register_inst104 <= 32'h0;	// <stdin>:5650:17, :5755:7
      Register_inst105 <= 32'h0;	// <stdin>:5650:17, :5756:7
      Register_inst106 <= 32'h0;	// <stdin>:5650:17, :5757:7
      Register_inst107 <= 32'h0;	// <stdin>:5650:17, :5758:7
      Register_inst108 <= 32'h0;	// <stdin>:5650:17, :5759:7
      Register_inst109 <= 32'h0;	// <stdin>:5650:17, :5760:7
      Register_inst110 <= 32'h0;	// <stdin>:5650:17, :5761:7
      Register_inst111 <= 32'h0;	// <stdin>:5650:17, :5762:7
      Register_inst112 <= 32'h0;	// <stdin>:5650:17, :5763:7
      Register_inst113 <= 32'h0;	// <stdin>:5650:17, :5764:7
      Register_inst114 <= 32'h0;	// <stdin>:5650:17, :5765:7
      Register_inst115 <= 32'h0;	// <stdin>:5650:17, :5766:7
      Register_inst116 <= 32'h0;	// <stdin>:5650:17, :5767:7
      Register_inst117 <= 32'h0;	// <stdin>:5650:17, :5768:7
      Register_inst118 <= 32'h0;	// <stdin>:5650:17, :5769:7
      Register_inst119 <= 32'h0;	// <stdin>:5650:17, :5770:7
      Register_inst120 <= 32'h0;	// <stdin>:5650:17, :5771:7
      Register_inst121 <= 32'h0;	// <stdin>:5650:17, :5772:7
      Register_inst122 <= 32'h0;	// <stdin>:5650:17, :5773:7
      Register_inst123 <= 32'h0;	// <stdin>:5650:17, :5774:7
      Register_inst124 <= 32'h0;	// <stdin>:5650:17, :5775:7
      Register_inst125 <= 32'h0;	// <stdin>:5650:17, :5776:7
      Register_inst126 <= 32'h0;	// <stdin>:5650:17, :5777:7
      Register_inst127 <= 32'h0;	// <stdin>:5650:17, :5778:7
      Register_inst128 <= 32'h0;	// <stdin>:5650:17, :5779:7
      Register_inst129 <= 32'h0;	// <stdin>:5650:17, :5780:7
      Register_inst130 <= 32'h0;	// <stdin>:5650:17, :5781:7
      Register_inst131 <= 32'h0;	// <stdin>:5650:17, :5782:7
      Register_inst132 <= 32'h0;	// <stdin>:5650:17, :5783:7
      Register_inst133 <= 32'h0;	// <stdin>:5650:17, :5784:7
      Register_inst134 <= 32'h0;	// <stdin>:5650:17, :5785:7
      Register_inst135 <= 32'h0;	// <stdin>:5650:17, :5786:7
      Register_inst136 <= 32'h0;	// <stdin>:5650:17, :5787:7
      Register_inst137 <= 32'h0;	// <stdin>:5650:17, :5788:7
      Register_inst138 <= 32'h0;	// <stdin>:5650:17, :5789:7
      Register_inst139 <= 32'h0;	// <stdin>:5650:17, :5790:7
      Register_inst140 <= 32'h0;	// <stdin>:5650:17, :5791:7
      Register_inst141 <= 32'h0;	// <stdin>:5650:17, :5792:7
      Register_inst142 <= 32'h0;	// <stdin>:5650:17, :5793:7
      Register_inst143 <= 32'h0;	// <stdin>:5650:17, :5794:7
      Register_inst144 <= 32'h0;	// <stdin>:5650:17, :5795:7
      Register_inst145 <= 32'h0;	// <stdin>:5650:17, :5796:7
      Register_inst146 <= 32'h0;	// <stdin>:5650:17, :5797:7
      Register_inst147 <= 32'h0;	// <stdin>:5650:17, :5798:7
      Register_inst148 <= 32'h0;	// <stdin>:5650:17, :5799:7
      Register_inst149 <= 32'h0;	// <stdin>:5650:17, :5800:7
      Register_inst150 <= 32'h0;	// <stdin>:5650:17, :5801:7
      Register_inst151 <= 32'h0;	// <stdin>:5650:17, :5802:7
      Register_inst152 <= 32'h0;	// <stdin>:5650:17, :5803:7
      Register_inst153 <= 32'h0;	// <stdin>:5650:17, :5804:7
      Register_inst154 <= 32'h0;	// <stdin>:5650:17, :5805:7
      Register_inst155 <= 32'h0;	// <stdin>:5650:17, :5806:7
      Register_inst156 <= 32'h0;	// <stdin>:5650:17, :5807:7
      Register_inst157 <= 32'h0;	// <stdin>:5650:17, :5808:7
      Register_inst158 <= 32'h0;	// <stdin>:5650:17, :5809:7
      Register_inst159 <= 32'h0;	// <stdin>:5650:17, :5810:7
      Register_inst160 <= 32'h0;	// <stdin>:5650:17, :5811:7
      Register_inst161 <= 32'h0;	// <stdin>:5650:17, :5812:7
      Register_inst162 <= 32'h0;	// <stdin>:5650:17, :5813:7
      Register_inst163 <= 32'h0;	// <stdin>:5650:17, :5814:7
      Register_inst164 <= 32'h0;	// <stdin>:5650:17, :5815:7
      Register_inst165 <= 32'h0;	// <stdin>:5650:17, :5816:7
      Register_inst166 <= 32'h0;	// <stdin>:5650:17, :5817:7
      Register_inst167 <= 32'h0;	// <stdin>:5650:17, :5818:7
      Register_inst168 <= 32'h0;	// <stdin>:5650:17, :5819:7
      Register_inst169 <= 32'h0;	// <stdin>:5650:17, :5820:7
      Register_inst170 <= 32'h0;	// <stdin>:5650:17, :5821:7
      Register_inst171 <= 32'h0;	// <stdin>:5650:17, :5822:7
      Register_inst172 <= 32'h0;	// <stdin>:5650:17, :5823:7
      Register_inst173 <= 32'h0;	// <stdin>:5650:17, :5824:7
      Register_inst174 <= 32'h0;	// <stdin>:5650:17, :5825:7
      Register_inst175 <= 32'h0;	// <stdin>:5650:17, :5826:7
      Register_inst176 <= 32'h0;	// <stdin>:5650:17, :5827:7
      Register_inst177 <= 32'h0;	// <stdin>:5650:17, :5828:7
      Register_inst178 <= 32'h0;	// <stdin>:5650:17, :5829:7
      Register_inst179 <= 32'h0;	// <stdin>:5650:17, :5830:7
      Register_inst180 <= 32'h0;	// <stdin>:5650:17, :5831:7
      Register_inst181 <= 32'h0;	// <stdin>:5650:17, :5832:7
      Register_inst182 <= 32'h0;	// <stdin>:5650:17, :5833:7
      Register_inst183 <= 32'h0;	// <stdin>:5650:17, :5834:7
      Register_inst184 <= 32'h0;	// <stdin>:5650:17, :5835:7
      Register_inst185 <= 32'h0;	// <stdin>:5650:17, :5836:7
      Register_inst186 <= 32'h0;	// <stdin>:5650:17, :5837:7
      Register_inst187 <= 32'h0;	// <stdin>:5650:17, :5838:7
      Register_inst188 <= 32'h0;	// <stdin>:5650:17, :5839:7
      Register_inst189 <= 32'h0;	// <stdin>:5650:17, :5840:7
      Register_inst190 <= 32'h0;	// <stdin>:5650:17, :5841:7
      Register_inst191 <= 32'h0;	// <stdin>:5650:17, :5842:7
      Register_inst192 <= 32'h0;	// <stdin>:5650:17, :5843:7
      Register_inst193 <= 32'h0;	// <stdin>:5650:17, :5844:7
      Register_inst194 <= 32'h0;	// <stdin>:5650:17, :5845:7
      Register_inst195 <= 32'h0;	// <stdin>:5650:17, :5846:7
      Register_inst196 <= 32'h0;	// <stdin>:5650:17, :5847:7
      Register_inst197 <= 32'h0;	// <stdin>:5650:17, :5848:7
      Register_inst198 <= 32'h0;	// <stdin>:5650:17, :5849:7
      Register_inst199 <= 32'h0;	// <stdin>:5650:17, :5850:7
      Register_inst200 <= 32'h0;	// <stdin>:5650:17, :5851:7
      Register_inst201 <= 32'h0;	// <stdin>:5650:17, :5852:7
      Register_inst202 <= 32'h0;	// <stdin>:5650:17, :5853:7
      Register_inst203 <= 32'h0;	// <stdin>:5650:17, :5854:7
      Register_inst204 <= 32'h0;	// <stdin>:5650:17, :5855:7
      Register_inst205 <= 32'h0;	// <stdin>:5650:17, :5856:7
      Register_inst206 <= 32'h0;	// <stdin>:5650:17, :5857:7
      Register_inst207 <= 32'h0;	// <stdin>:5650:17, :5858:7
      Register_inst208 <= 32'h0;	// <stdin>:5650:17, :5859:7
      Register_inst209 <= 32'h0;	// <stdin>:5650:17, :5860:7
      Register_inst210 <= 32'h0;	// <stdin>:5650:17, :5861:7
      Register_inst211 <= 32'h0;	// <stdin>:5650:17, :5862:7
      Register_inst212 <= 32'h0;	// <stdin>:5650:17, :5863:7
      Register_inst213 <= 32'h0;	// <stdin>:5650:17, :5864:7
      Register_inst214 <= 32'h0;	// <stdin>:5650:17, :5865:7
      Register_inst215 <= 32'h0;	// <stdin>:5650:17, :5866:7
      Register_inst216 <= 32'h0;	// <stdin>:5650:17, :5867:7
      Register_inst217 <= 32'h0;	// <stdin>:5650:17, :5868:7
      Register_inst218 <= 32'h0;	// <stdin>:5650:17, :5869:7
      Register_inst219 <= 32'h0;	// <stdin>:5650:17, :5870:7
      Register_inst220 <= 32'h0;	// <stdin>:5650:17, :5871:7
      Register_inst221 <= 32'h0;	// <stdin>:5650:17, :5872:7
      Register_inst222 <= 32'h0;	// <stdin>:5650:17, :5873:7
      Register_inst223 <= 32'h0;	// <stdin>:5650:17, :5874:7
      Register_inst224 <= 32'h0;	// <stdin>:5650:17, :5875:7
      Register_inst225 <= 32'h0;	// <stdin>:5650:17, :5876:7
      Register_inst226 <= 32'h0;	// <stdin>:5650:17, :5877:7
      Register_inst227 <= 32'h0;	// <stdin>:5650:17, :5878:7
      Register_inst228 <= 32'h0;	// <stdin>:5650:17, :5879:7
      Register_inst229 <= 32'h0;	// <stdin>:5650:17, :5880:7
      Register_inst230 <= 32'h0;	// <stdin>:5650:17, :5881:7
      Register_inst231 <= 32'h0;	// <stdin>:5650:17, :5882:7
      Register_inst232 <= 32'h0;	// <stdin>:5650:17, :5883:7
      Register_inst233 <= 32'h0;	// <stdin>:5650:17, :5884:7
      Register_inst234 <= 32'h0;	// <stdin>:5650:17, :5885:7
      Register_inst235 <= 32'h0;	// <stdin>:5650:17, :5886:7
      Register_inst236 <= 32'h0;	// <stdin>:5650:17, :5887:7
      Register_inst237 <= 32'h0;	// <stdin>:5650:17, :5888:7
      Register_inst238 <= 32'h0;	// <stdin>:5650:17, :5889:7
      Register_inst239 <= 32'h0;	// <stdin>:5650:17, :5890:7
      Register_inst240 <= 32'h0;	// <stdin>:5650:17, :5891:7
      Register_inst241 <= 32'h0;	// <stdin>:5650:17, :5892:7
      Register_inst242 <= 32'h0;	// <stdin>:5650:17, :5893:7
      Register_inst243 <= 32'h0;	// <stdin>:5650:17, :5894:7
      Register_inst244 <= 32'h0;	// <stdin>:5650:17, :5895:7
      Register_inst245 <= 32'h0;	// <stdin>:5650:17, :5896:7
      Register_inst246 <= 32'h0;	// <stdin>:5650:17, :5897:7
      Register_inst247 <= 32'h0;	// <stdin>:5650:17, :5898:7
      Register_inst248 <= 32'h0;	// <stdin>:5650:17, :5899:7
      Register_inst249 <= 32'h0;	// <stdin>:5650:17, :5900:7
      Register_inst250 <= 32'h0;	// <stdin>:5650:17, :5901:7
      Register_inst251 <= 32'h0;	// <stdin>:5650:17, :5902:7
      Register_inst252 <= 32'h0;	// <stdin>:5650:17, :5903:7
      Register_inst253 <= 32'h0;	// <stdin>:5650:17, :5904:7
      Register_inst254 <= 32'h0;	// <stdin>:5650:17, :5905:7
      Register_inst255 <= 32'h0;	// <stdin>:5650:17, :5906:7
    end
    else begin	// <stdin>:5392:5
      Register_inst0 <= _T_255;	// <stdin>:5393:7
      Register_inst1 <= _T_256;	// <stdin>:5394:7
      Register_inst2 <= _T_257;	// <stdin>:5395:7
      Register_inst3 <= _T_258;	// <stdin>:5396:7
      Register_inst4 <= _T_259;	// <stdin>:5397:7
      Register_inst5 <= _T_260;	// <stdin>:5398:7
      Register_inst6 <= _T_261;	// <stdin>:5399:7
      Register_inst7 <= _T_262;	// <stdin>:5400:7
      Register_inst8 <= _T_263;	// <stdin>:5401:7
      Register_inst9 <= _T_264;	// <stdin>:5402:7
      Register_inst10 <= _T_265;	// <stdin>:5403:7
      Register_inst11 <= _T_266;	// <stdin>:5404:7
      Register_inst12 <= _T_267;	// <stdin>:5405:7
      Register_inst13 <= _T_268;	// <stdin>:5406:7
      Register_inst14 <= _T_269;	// <stdin>:5407:7
      Register_inst15 <= _T_270;	// <stdin>:5408:7
      Register_inst16 <= _T_271;	// <stdin>:5409:7
      Register_inst17 <= _T_272;	// <stdin>:5410:7
      Register_inst18 <= _T_273;	// <stdin>:5411:7
      Register_inst19 <= _T_274;	// <stdin>:5412:7
      Register_inst20 <= _T_275;	// <stdin>:5413:7
      Register_inst21 <= _T_276;	// <stdin>:5414:7
      Register_inst22 <= _T_277;	// <stdin>:5415:7
      Register_inst23 <= _T_278;	// <stdin>:5416:7
      Register_inst24 <= _T_279;	// <stdin>:5417:7
      Register_inst25 <= _T_280;	// <stdin>:5418:7
      Register_inst26 <= _T_281;	// <stdin>:5419:7
      Register_inst27 <= _T_282;	// <stdin>:5420:7
      Register_inst28 <= _T_283;	// <stdin>:5421:7
      Register_inst29 <= _T_284;	// <stdin>:5422:7
      Register_inst30 <= _T_285;	// <stdin>:5423:7
      Register_inst31 <= _T_286;	// <stdin>:5424:7
      Register_inst32 <= _T_287;	// <stdin>:5425:7
      Register_inst33 <= _T_288;	// <stdin>:5426:7
      Register_inst34 <= _T_289;	// <stdin>:5427:7
      Register_inst35 <= _T_290;	// <stdin>:5428:7
      Register_inst36 <= _T_291;	// <stdin>:5429:7
      Register_inst37 <= _T_292;	// <stdin>:5430:7
      Register_inst38 <= _T_293;	// <stdin>:5431:7
      Register_inst39 <= _T_294;	// <stdin>:5432:7
      Register_inst40 <= _T_295;	// <stdin>:5433:7
      Register_inst41 <= _T_296;	// <stdin>:5434:7
      Register_inst42 <= _T_297;	// <stdin>:5435:7
      Register_inst43 <= _T_298;	// <stdin>:5436:7
      Register_inst44 <= _T_299;	// <stdin>:5437:7
      Register_inst45 <= _T_300;	// <stdin>:5438:7
      Register_inst46 <= _T_301;	// <stdin>:5439:7
      Register_inst47 <= _T_302;	// <stdin>:5440:7
      Register_inst48 <= _T_303;	// <stdin>:5441:7
      Register_inst49 <= _T_304;	// <stdin>:5442:7
      Register_inst50 <= _T_305;	// <stdin>:5443:7
      Register_inst51 <= _T_306;	// <stdin>:5444:7
      Register_inst52 <= _T_307;	// <stdin>:5445:7
      Register_inst53 <= _T_308;	// <stdin>:5446:7
      Register_inst54 <= _T_309;	// <stdin>:5447:7
      Register_inst55 <= _T_310;	// <stdin>:5448:7
      Register_inst56 <= _T_311;	// <stdin>:5449:7
      Register_inst57 <= _T_312;	// <stdin>:5450:7
      Register_inst58 <= _T_313;	// <stdin>:5451:7
      Register_inst59 <= _T_314;	// <stdin>:5452:7
      Register_inst60 <= _T_315;	// <stdin>:5453:7
      Register_inst61 <= _T_316;	// <stdin>:5454:7
      Register_inst62 <= _T_317;	// <stdin>:5455:7
      Register_inst63 <= _T_318;	// <stdin>:5456:7
      Register_inst64 <= _T_319;	// <stdin>:5457:7
      Register_inst65 <= _T_320;	// <stdin>:5458:7
      Register_inst66 <= _T_321;	// <stdin>:5459:7
      Register_inst67 <= _T_322;	// <stdin>:5460:7
      Register_inst68 <= _T_323;	// <stdin>:5461:7
      Register_inst69 <= _T_324;	// <stdin>:5462:7
      Register_inst70 <= _T_325;	// <stdin>:5463:7
      Register_inst71 <= _T_326;	// <stdin>:5464:7
      Register_inst72 <= _T_327;	// <stdin>:5465:7
      Register_inst73 <= _T_328;	// <stdin>:5466:7
      Register_inst74 <= _T_329;	// <stdin>:5467:7
      Register_inst75 <= _T_330;	// <stdin>:5468:7
      Register_inst76 <= _T_331;	// <stdin>:5469:7
      Register_inst77 <= _T_332;	// <stdin>:5470:7
      Register_inst78 <= _T_333;	// <stdin>:5471:7
      Register_inst79 <= _T_334;	// <stdin>:5472:7
      Register_inst80 <= _T_335;	// <stdin>:5473:7
      Register_inst81 <= _T_336;	// <stdin>:5474:7
      Register_inst82 <= _T_337;	// <stdin>:5475:7
      Register_inst83 <= _T_338;	// <stdin>:5476:7
      Register_inst84 <= _T_339;	// <stdin>:5477:7
      Register_inst85 <= _T_340;	// <stdin>:5478:7
      Register_inst86 <= _T_341;	// <stdin>:5479:7
      Register_inst87 <= _T_342;	// <stdin>:5480:7
      Register_inst88 <= _T_343;	// <stdin>:5481:7
      Register_inst89 <= _T_344;	// <stdin>:5482:7
      Register_inst90 <= _T_345;	// <stdin>:5483:7
      Register_inst91 <= _T_346;	// <stdin>:5484:7
      Register_inst92 <= _T_347;	// <stdin>:5485:7
      Register_inst93 <= _T_348;	// <stdin>:5486:7
      Register_inst94 <= _T_349;	// <stdin>:5487:7
      Register_inst95 <= _T_350;	// <stdin>:5488:7
      Register_inst96 <= _T_351;	// <stdin>:5489:7
      Register_inst97 <= _T_352;	// <stdin>:5490:7
      Register_inst98 <= _T_353;	// <stdin>:5491:7
      Register_inst99 <= _T_354;	// <stdin>:5492:7
      Register_inst100 <= _T_355;	// <stdin>:5493:7
      Register_inst101 <= _T_356;	// <stdin>:5494:7
      Register_inst102 <= _T_357;	// <stdin>:5495:7
      Register_inst103 <= _T_358;	// <stdin>:5496:7
      Register_inst104 <= _T_359;	// <stdin>:5497:7
      Register_inst105 <= _T_360;	// <stdin>:5498:7
      Register_inst106 <= _T_361;	// <stdin>:5499:7
      Register_inst107 <= _T_362;	// <stdin>:5500:7
      Register_inst108 <= _T_363;	// <stdin>:5501:7
      Register_inst109 <= _T_364;	// <stdin>:5502:7
      Register_inst110 <= _T_365;	// <stdin>:5503:7
      Register_inst111 <= _T_366;	// <stdin>:5504:7
      Register_inst112 <= _T_367;	// <stdin>:5505:7
      Register_inst113 <= _T_368;	// <stdin>:5506:7
      Register_inst114 <= _T_369;	// <stdin>:5507:7
      Register_inst115 <= _T_370;	// <stdin>:5508:7
      Register_inst116 <= _T_371;	// <stdin>:5509:7
      Register_inst117 <= _T_372;	// <stdin>:5510:7
      Register_inst118 <= _T_373;	// <stdin>:5511:7
      Register_inst119 <= _T_374;	// <stdin>:5512:7
      Register_inst120 <= _T_375;	// <stdin>:5513:7
      Register_inst121 <= _T_376;	// <stdin>:5514:7
      Register_inst122 <= _T_377;	// <stdin>:5515:7
      Register_inst123 <= _T_378;	// <stdin>:5516:7
      Register_inst124 <= _T_379;	// <stdin>:5517:7
      Register_inst125 <= _T_380;	// <stdin>:5518:7
      Register_inst126 <= _T_381;	// <stdin>:5519:7
      Register_inst127 <= _T_382;	// <stdin>:5520:7
      Register_inst128 <= _T_383;	// <stdin>:5521:7
      Register_inst129 <= _T_384;	// <stdin>:5522:7
      Register_inst130 <= _T_385;	// <stdin>:5523:7
      Register_inst131 <= _T_386;	// <stdin>:5524:7
      Register_inst132 <= _T_387;	// <stdin>:5525:7
      Register_inst133 <= _T_388;	// <stdin>:5526:7
      Register_inst134 <= _T_389;	// <stdin>:5527:7
      Register_inst135 <= _T_390;	// <stdin>:5528:7
      Register_inst136 <= _T_391;	// <stdin>:5529:7
      Register_inst137 <= _T_392;	// <stdin>:5530:7
      Register_inst138 <= _T_393;	// <stdin>:5531:7
      Register_inst139 <= _T_394;	// <stdin>:5532:7
      Register_inst140 <= _T_395;	// <stdin>:5533:7
      Register_inst141 <= _T_396;	// <stdin>:5534:7
      Register_inst142 <= _T_397;	// <stdin>:5535:7
      Register_inst143 <= _T_398;	// <stdin>:5536:7
      Register_inst144 <= _T_399;	// <stdin>:5537:7
      Register_inst145 <= _T_400;	// <stdin>:5538:7
      Register_inst146 <= _T_401;	// <stdin>:5539:7
      Register_inst147 <= _T_402;	// <stdin>:5540:7
      Register_inst148 <= _T_403;	// <stdin>:5541:7
      Register_inst149 <= _T_404;	// <stdin>:5542:7
      Register_inst150 <= _T_405;	// <stdin>:5543:7
      Register_inst151 <= _T_406;	// <stdin>:5544:7
      Register_inst152 <= _T_407;	// <stdin>:5545:7
      Register_inst153 <= _T_408;	// <stdin>:5546:7
      Register_inst154 <= _T_409;	// <stdin>:5547:7
      Register_inst155 <= _T_410;	// <stdin>:5548:7
      Register_inst156 <= _T_411;	// <stdin>:5549:7
      Register_inst157 <= _T_412;	// <stdin>:5550:7
      Register_inst158 <= _T_413;	// <stdin>:5551:7
      Register_inst159 <= _T_414;	// <stdin>:5552:7
      Register_inst160 <= _T_415;	// <stdin>:5553:7
      Register_inst161 <= _T_416;	// <stdin>:5554:7
      Register_inst162 <= _T_417;	// <stdin>:5555:7
      Register_inst163 <= _T_418;	// <stdin>:5556:7
      Register_inst164 <= _T_419;	// <stdin>:5557:7
      Register_inst165 <= _T_420;	// <stdin>:5558:7
      Register_inst166 <= _T_421;	// <stdin>:5559:7
      Register_inst167 <= _T_422;	// <stdin>:5560:7
      Register_inst168 <= _T_423;	// <stdin>:5561:7
      Register_inst169 <= _T_424;	// <stdin>:5562:7
      Register_inst170 <= _T_425;	// <stdin>:5563:7
      Register_inst171 <= _T_426;	// <stdin>:5564:7
      Register_inst172 <= _T_427;	// <stdin>:5565:7
      Register_inst173 <= _T_428;	// <stdin>:5566:7
      Register_inst174 <= _T_429;	// <stdin>:5567:7
      Register_inst175 <= _T_430;	// <stdin>:5568:7
      Register_inst176 <= _T_431;	// <stdin>:5569:7
      Register_inst177 <= _T_432;	// <stdin>:5570:7
      Register_inst178 <= _T_433;	// <stdin>:5571:7
      Register_inst179 <= _T_434;	// <stdin>:5572:7
      Register_inst180 <= _T_435;	// <stdin>:5573:7
      Register_inst181 <= _T_436;	// <stdin>:5574:7
      Register_inst182 <= _T_437;	// <stdin>:5575:7
      Register_inst183 <= _T_438;	// <stdin>:5576:7
      Register_inst184 <= _T_439;	// <stdin>:5577:7
      Register_inst185 <= _T_440;	// <stdin>:5578:7
      Register_inst186 <= _T_441;	// <stdin>:5579:7
      Register_inst187 <= _T_442;	// <stdin>:5580:7
      Register_inst188 <= _T_443;	// <stdin>:5581:7
      Register_inst189 <= _T_444;	// <stdin>:5582:7
      Register_inst190 <= _T_445;	// <stdin>:5583:7
      Register_inst191 <= _T_446;	// <stdin>:5584:7
      Register_inst192 <= _T_447;	// <stdin>:5585:7
      Register_inst193 <= _T_448;	// <stdin>:5586:7
      Register_inst194 <= _T_449;	// <stdin>:5587:7
      Register_inst195 <= _T_450;	// <stdin>:5588:7
      Register_inst196 <= _T_451;	// <stdin>:5589:7
      Register_inst197 <= _T_452;	// <stdin>:5590:7
      Register_inst198 <= _T_453;	// <stdin>:5591:7
      Register_inst199 <= _T_454;	// <stdin>:5592:7
      Register_inst200 <= _T_455;	// <stdin>:5593:7
      Register_inst201 <= _T_456;	// <stdin>:5594:7
      Register_inst202 <= _T_457;	// <stdin>:5595:7
      Register_inst203 <= _T_458;	// <stdin>:5596:7
      Register_inst204 <= _T_459;	// <stdin>:5597:7
      Register_inst205 <= _T_460;	// <stdin>:5598:7
      Register_inst206 <= _T_461;	// <stdin>:5599:7
      Register_inst207 <= _T_462;	// <stdin>:5600:7
      Register_inst208 <= _T_463;	// <stdin>:5601:7
      Register_inst209 <= _T_464;	// <stdin>:5602:7
      Register_inst210 <= _T_465;	// <stdin>:5603:7
      Register_inst211 <= _T_466;	// <stdin>:5604:7
      Register_inst212 <= _T_467;	// <stdin>:5605:7
      Register_inst213 <= _T_468;	// <stdin>:5606:7
      Register_inst214 <= _T_469;	// <stdin>:5607:7
      Register_inst215 <= _T_470;	// <stdin>:5608:7
      Register_inst216 <= _T_471;	// <stdin>:5609:7
      Register_inst217 <= _T_472;	// <stdin>:5610:7
      Register_inst218 <= _T_473;	// <stdin>:5611:7
      Register_inst219 <= _T_474;	// <stdin>:5612:7
      Register_inst220 <= _T_475;	// <stdin>:5613:7
      Register_inst221 <= _T_476;	// <stdin>:5614:7
      Register_inst222 <= _T_477;	// <stdin>:5615:7
      Register_inst223 <= _T_478;	// <stdin>:5616:7
      Register_inst224 <= _T_479;	// <stdin>:5617:7
      Register_inst225 <= _T_480;	// <stdin>:5618:7
      Register_inst226 <= _T_481;	// <stdin>:5619:7
      Register_inst227 <= _T_482;	// <stdin>:5620:7
      Register_inst228 <= _T_483;	// <stdin>:5621:7
      Register_inst229 <= _T_484;	// <stdin>:5622:7
      Register_inst230 <= _T_485;	// <stdin>:5623:7
      Register_inst231 <= _T_486;	// <stdin>:5624:7
      Register_inst232 <= _T_487;	// <stdin>:5625:7
      Register_inst233 <= _T_488;	// <stdin>:5626:7
      Register_inst234 <= _T_489;	// <stdin>:5627:7
      Register_inst235 <= _T_490;	// <stdin>:5628:7
      Register_inst236 <= _T_491;	// <stdin>:5629:7
      Register_inst237 <= _T_492;	// <stdin>:5630:7
      Register_inst238 <= _T_493;	// <stdin>:5631:7
      Register_inst239 <= _T_494;	// <stdin>:5632:7
      Register_inst240 <= _T_495;	// <stdin>:5633:7
      Register_inst241 <= _T_496;	// <stdin>:5634:7
      Register_inst242 <= _T_497;	// <stdin>:5635:7
      Register_inst243 <= _T_498;	// <stdin>:5636:7
      Register_inst244 <= _T_499;	// <stdin>:5637:7
      Register_inst245 <= _T_500;	// <stdin>:5638:7
      Register_inst246 <= _T_501;	// <stdin>:5639:7
      Register_inst247 <= _T_502;	// <stdin>:5640:7
      Register_inst248 <= _T_503;	// <stdin>:5641:7
      Register_inst249 <= _T_504;	// <stdin>:5642:7
      Register_inst250 <= _T_505;	// <stdin>:5643:7
      Register_inst251 <= _T_506;	// <stdin>:5644:7
      Register_inst252 <= _T_507;	// <stdin>:5645:7
      Register_inst253 <= _T_508;	// <stdin>:5646:7
      Register_inst254 <= _T_509;	// <stdin>:5647:7
      Register_inst255 <= _T_510;	// <stdin>:5648:7
    end
  end // always @(posedge or posedge)
  initial begin	// <stdin>:5908:5
    Register_inst0 = 32'h0;	// <stdin>:5909:17, :5910:7
    Register_inst1 = 32'h0;	// <stdin>:5909:17, :5911:7
    Register_inst2 = 32'h0;	// <stdin>:5909:17, :5912:7
    Register_inst3 = 32'h0;	// <stdin>:5909:17, :5913:7
    Register_inst4 = 32'h0;	// <stdin>:5909:17, :5914:7
    Register_inst5 = 32'h0;	// <stdin>:5909:17, :5915:7
    Register_inst6 = 32'h0;	// <stdin>:5909:17, :5916:7
    Register_inst7 = 32'h0;	// <stdin>:5909:17, :5917:7
    Register_inst8 = 32'h0;	// <stdin>:5909:17, :5918:7
    Register_inst9 = 32'h0;	// <stdin>:5909:17, :5919:7
    Register_inst10 = 32'h0;	// <stdin>:5909:17, :5920:7
    Register_inst11 = 32'h0;	// <stdin>:5909:17, :5921:7
    Register_inst12 = 32'h0;	// <stdin>:5909:17, :5922:7
    Register_inst13 = 32'h0;	// <stdin>:5909:17, :5923:7
    Register_inst14 = 32'h0;	// <stdin>:5909:17, :5924:7
    Register_inst15 = 32'h0;	// <stdin>:5909:17, :5925:7
    Register_inst16 = 32'h0;	// <stdin>:5909:17, :5926:7
    Register_inst17 = 32'h0;	// <stdin>:5909:17, :5927:7
    Register_inst18 = 32'h0;	// <stdin>:5909:17, :5928:7
    Register_inst19 = 32'h0;	// <stdin>:5909:17, :5929:7
    Register_inst20 = 32'h0;	// <stdin>:5909:17, :5930:7
    Register_inst21 = 32'h0;	// <stdin>:5909:17, :5931:7
    Register_inst22 = 32'h0;	// <stdin>:5909:17, :5932:7
    Register_inst23 = 32'h0;	// <stdin>:5909:17, :5933:7
    Register_inst24 = 32'h0;	// <stdin>:5909:17, :5934:7
    Register_inst25 = 32'h0;	// <stdin>:5909:17, :5935:7
    Register_inst26 = 32'h0;	// <stdin>:5909:17, :5936:7
    Register_inst27 = 32'h0;	// <stdin>:5909:17, :5937:7
    Register_inst28 = 32'h0;	// <stdin>:5909:17, :5938:7
    Register_inst29 = 32'h0;	// <stdin>:5909:17, :5939:7
    Register_inst30 = 32'h0;	// <stdin>:5909:17, :5940:7
    Register_inst31 = 32'h0;	// <stdin>:5909:17, :5941:7
    Register_inst32 = 32'h0;	// <stdin>:5909:17, :5942:7
    Register_inst33 = 32'h0;	// <stdin>:5909:17, :5943:7
    Register_inst34 = 32'h0;	// <stdin>:5909:17, :5944:7
    Register_inst35 = 32'h0;	// <stdin>:5909:17, :5945:7
    Register_inst36 = 32'h0;	// <stdin>:5909:17, :5946:7
    Register_inst37 = 32'h0;	// <stdin>:5909:17, :5947:7
    Register_inst38 = 32'h0;	// <stdin>:5909:17, :5948:7
    Register_inst39 = 32'h0;	// <stdin>:5909:17, :5949:7
    Register_inst40 = 32'h0;	// <stdin>:5909:17, :5950:7
    Register_inst41 = 32'h0;	// <stdin>:5909:17, :5951:7
    Register_inst42 = 32'h0;	// <stdin>:5909:17, :5952:7
    Register_inst43 = 32'h0;	// <stdin>:5909:17, :5953:7
    Register_inst44 = 32'h0;	// <stdin>:5909:17, :5954:7
    Register_inst45 = 32'h0;	// <stdin>:5909:17, :5955:7
    Register_inst46 = 32'h0;	// <stdin>:5909:17, :5956:7
    Register_inst47 = 32'h0;	// <stdin>:5909:17, :5957:7
    Register_inst48 = 32'h0;	// <stdin>:5909:17, :5958:7
    Register_inst49 = 32'h0;	// <stdin>:5909:17, :5959:7
    Register_inst50 = 32'h0;	// <stdin>:5909:17, :5960:7
    Register_inst51 = 32'h0;	// <stdin>:5909:17, :5961:7
    Register_inst52 = 32'h0;	// <stdin>:5909:17, :5962:7
    Register_inst53 = 32'h0;	// <stdin>:5909:17, :5963:7
    Register_inst54 = 32'h0;	// <stdin>:5909:17, :5964:7
    Register_inst55 = 32'h0;	// <stdin>:5909:17, :5965:7
    Register_inst56 = 32'h0;	// <stdin>:5909:17, :5966:7
    Register_inst57 = 32'h0;	// <stdin>:5909:17, :5967:7
    Register_inst58 = 32'h0;	// <stdin>:5909:17, :5968:7
    Register_inst59 = 32'h0;	// <stdin>:5909:17, :5969:7
    Register_inst60 = 32'h0;	// <stdin>:5909:17, :5970:7
    Register_inst61 = 32'h0;	// <stdin>:5909:17, :5971:7
    Register_inst62 = 32'h0;	// <stdin>:5909:17, :5972:7
    Register_inst63 = 32'h0;	// <stdin>:5909:17, :5973:7
    Register_inst64 = 32'h0;	// <stdin>:5909:17, :5974:7
    Register_inst65 = 32'h0;	// <stdin>:5909:17, :5975:7
    Register_inst66 = 32'h0;	// <stdin>:5909:17, :5976:7
    Register_inst67 = 32'h0;	// <stdin>:5909:17, :5977:7
    Register_inst68 = 32'h0;	// <stdin>:5909:17, :5978:7
    Register_inst69 = 32'h0;	// <stdin>:5909:17, :5979:7
    Register_inst70 = 32'h0;	// <stdin>:5909:17, :5980:7
    Register_inst71 = 32'h0;	// <stdin>:5909:17, :5981:7
    Register_inst72 = 32'h0;	// <stdin>:5909:17, :5982:7
    Register_inst73 = 32'h0;	// <stdin>:5909:17, :5983:7
    Register_inst74 = 32'h0;	// <stdin>:5909:17, :5984:7
    Register_inst75 = 32'h0;	// <stdin>:5909:17, :5985:7
    Register_inst76 = 32'h0;	// <stdin>:5909:17, :5986:7
    Register_inst77 = 32'h0;	// <stdin>:5909:17, :5987:7
    Register_inst78 = 32'h0;	// <stdin>:5909:17, :5988:7
    Register_inst79 = 32'h0;	// <stdin>:5909:17, :5989:7
    Register_inst80 = 32'h0;	// <stdin>:5909:17, :5990:7
    Register_inst81 = 32'h0;	// <stdin>:5909:17, :5991:7
    Register_inst82 = 32'h0;	// <stdin>:5909:17, :5992:7
    Register_inst83 = 32'h0;	// <stdin>:5909:17, :5993:7
    Register_inst84 = 32'h0;	// <stdin>:5909:17, :5994:7
    Register_inst85 = 32'h0;	// <stdin>:5909:17, :5995:7
    Register_inst86 = 32'h0;	// <stdin>:5909:17, :5996:7
    Register_inst87 = 32'h0;	// <stdin>:5909:17, :5997:7
    Register_inst88 = 32'h0;	// <stdin>:5909:17, :5998:7
    Register_inst89 = 32'h0;	// <stdin>:5909:17, :5999:7
    Register_inst90 = 32'h0;	// <stdin>:5909:17, :6000:7
    Register_inst91 = 32'h0;	// <stdin>:5909:17, :6001:7
    Register_inst92 = 32'h0;	// <stdin>:5909:17, :6002:7
    Register_inst93 = 32'h0;	// <stdin>:5909:17, :6003:7
    Register_inst94 = 32'h0;	// <stdin>:5909:17, :6004:7
    Register_inst95 = 32'h0;	// <stdin>:5909:17, :6005:7
    Register_inst96 = 32'h0;	// <stdin>:5909:17, :6006:7
    Register_inst97 = 32'h0;	// <stdin>:5909:17, :6007:7
    Register_inst98 = 32'h0;	// <stdin>:5909:17, :6008:7
    Register_inst99 = 32'h0;	// <stdin>:5909:17, :6009:7
    Register_inst100 = 32'h0;	// <stdin>:5909:17, :6010:7
    Register_inst101 = 32'h0;	// <stdin>:5909:17, :6011:7
    Register_inst102 = 32'h0;	// <stdin>:5909:17, :6012:7
    Register_inst103 = 32'h0;	// <stdin>:5909:17, :6013:7
    Register_inst104 = 32'h0;	// <stdin>:5909:17, :6014:7
    Register_inst105 = 32'h0;	// <stdin>:5909:17, :6015:7
    Register_inst106 = 32'h0;	// <stdin>:5909:17, :6016:7
    Register_inst107 = 32'h0;	// <stdin>:5909:17, :6017:7
    Register_inst108 = 32'h0;	// <stdin>:5909:17, :6018:7
    Register_inst109 = 32'h0;	// <stdin>:5909:17, :6019:7
    Register_inst110 = 32'h0;	// <stdin>:5909:17, :6020:7
    Register_inst111 = 32'h0;	// <stdin>:5909:17, :6021:7
    Register_inst112 = 32'h0;	// <stdin>:5909:17, :6022:7
    Register_inst113 = 32'h0;	// <stdin>:5909:17, :6023:7
    Register_inst114 = 32'h0;	// <stdin>:5909:17, :6024:7
    Register_inst115 = 32'h0;	// <stdin>:5909:17, :6025:7
    Register_inst116 = 32'h0;	// <stdin>:5909:17, :6026:7
    Register_inst117 = 32'h0;	// <stdin>:5909:17, :6027:7
    Register_inst118 = 32'h0;	// <stdin>:5909:17, :6028:7
    Register_inst119 = 32'h0;	// <stdin>:5909:17, :6029:7
    Register_inst120 = 32'h0;	// <stdin>:5909:17, :6030:7
    Register_inst121 = 32'h0;	// <stdin>:5909:17, :6031:7
    Register_inst122 = 32'h0;	// <stdin>:5909:17, :6032:7
    Register_inst123 = 32'h0;	// <stdin>:5909:17, :6033:7
    Register_inst124 = 32'h0;	// <stdin>:5909:17, :6034:7
    Register_inst125 = 32'h0;	// <stdin>:5909:17, :6035:7
    Register_inst126 = 32'h0;	// <stdin>:5909:17, :6036:7
    Register_inst127 = 32'h0;	// <stdin>:5909:17, :6037:7
    Register_inst128 = 32'h0;	// <stdin>:5909:17, :6038:7
    Register_inst129 = 32'h0;	// <stdin>:5909:17, :6039:7
    Register_inst130 = 32'h0;	// <stdin>:5909:17, :6040:7
    Register_inst131 = 32'h0;	// <stdin>:5909:17, :6041:7
    Register_inst132 = 32'h0;	// <stdin>:5909:17, :6042:7
    Register_inst133 = 32'h0;	// <stdin>:5909:17, :6043:7
    Register_inst134 = 32'h0;	// <stdin>:5909:17, :6044:7
    Register_inst135 = 32'h0;	// <stdin>:5909:17, :6045:7
    Register_inst136 = 32'h0;	// <stdin>:5909:17, :6046:7
    Register_inst137 = 32'h0;	// <stdin>:5909:17, :6047:7
    Register_inst138 = 32'h0;	// <stdin>:5909:17, :6048:7
    Register_inst139 = 32'h0;	// <stdin>:5909:17, :6049:7
    Register_inst140 = 32'h0;	// <stdin>:5909:17, :6050:7
    Register_inst141 = 32'h0;	// <stdin>:5909:17, :6051:7
    Register_inst142 = 32'h0;	// <stdin>:5909:17, :6052:7
    Register_inst143 = 32'h0;	// <stdin>:5909:17, :6053:7
    Register_inst144 = 32'h0;	// <stdin>:5909:17, :6054:7
    Register_inst145 = 32'h0;	// <stdin>:5909:17, :6055:7
    Register_inst146 = 32'h0;	// <stdin>:5909:17, :6056:7
    Register_inst147 = 32'h0;	// <stdin>:5909:17, :6057:7
    Register_inst148 = 32'h0;	// <stdin>:5909:17, :6058:7
    Register_inst149 = 32'h0;	// <stdin>:5909:17, :6059:7
    Register_inst150 = 32'h0;	// <stdin>:5909:17, :6060:7
    Register_inst151 = 32'h0;	// <stdin>:5909:17, :6061:7
    Register_inst152 = 32'h0;	// <stdin>:5909:17, :6062:7
    Register_inst153 = 32'h0;	// <stdin>:5909:17, :6063:7
    Register_inst154 = 32'h0;	// <stdin>:5909:17, :6064:7
    Register_inst155 = 32'h0;	// <stdin>:5909:17, :6065:7
    Register_inst156 = 32'h0;	// <stdin>:5909:17, :6066:7
    Register_inst157 = 32'h0;	// <stdin>:5909:17, :6067:7
    Register_inst158 = 32'h0;	// <stdin>:5909:17, :6068:7
    Register_inst159 = 32'h0;	// <stdin>:5909:17, :6069:7
    Register_inst160 = 32'h0;	// <stdin>:5909:17, :6070:7
    Register_inst161 = 32'h0;	// <stdin>:5909:17, :6071:7
    Register_inst162 = 32'h0;	// <stdin>:5909:17, :6072:7
    Register_inst163 = 32'h0;	// <stdin>:5909:17, :6073:7
    Register_inst164 = 32'h0;	// <stdin>:5909:17, :6074:7
    Register_inst165 = 32'h0;	// <stdin>:5909:17, :6075:7
    Register_inst166 = 32'h0;	// <stdin>:5909:17, :6076:7
    Register_inst167 = 32'h0;	// <stdin>:5909:17, :6077:7
    Register_inst168 = 32'h0;	// <stdin>:5909:17, :6078:7
    Register_inst169 = 32'h0;	// <stdin>:5909:17, :6079:7
    Register_inst170 = 32'h0;	// <stdin>:5909:17, :6080:7
    Register_inst171 = 32'h0;	// <stdin>:5909:17, :6081:7
    Register_inst172 = 32'h0;	// <stdin>:5909:17, :6082:7
    Register_inst173 = 32'h0;	// <stdin>:5909:17, :6083:7
    Register_inst174 = 32'h0;	// <stdin>:5909:17, :6084:7
    Register_inst175 = 32'h0;	// <stdin>:5909:17, :6085:7
    Register_inst176 = 32'h0;	// <stdin>:5909:17, :6086:7
    Register_inst177 = 32'h0;	// <stdin>:5909:17, :6087:7
    Register_inst178 = 32'h0;	// <stdin>:5909:17, :6088:7
    Register_inst179 = 32'h0;	// <stdin>:5909:17, :6089:7
    Register_inst180 = 32'h0;	// <stdin>:5909:17, :6090:7
    Register_inst181 = 32'h0;	// <stdin>:5909:17, :6091:7
    Register_inst182 = 32'h0;	// <stdin>:5909:17, :6092:7
    Register_inst183 = 32'h0;	// <stdin>:5909:17, :6093:7
    Register_inst184 = 32'h0;	// <stdin>:5909:17, :6094:7
    Register_inst185 = 32'h0;	// <stdin>:5909:17, :6095:7
    Register_inst186 = 32'h0;	// <stdin>:5909:17, :6096:7
    Register_inst187 = 32'h0;	// <stdin>:5909:17, :6097:7
    Register_inst188 = 32'h0;	// <stdin>:5909:17, :6098:7
    Register_inst189 = 32'h0;	// <stdin>:5909:17, :6099:7
    Register_inst190 = 32'h0;	// <stdin>:5909:17, :6100:7
    Register_inst191 = 32'h0;	// <stdin>:5909:17, :6101:7
    Register_inst192 = 32'h0;	// <stdin>:5909:17, :6102:7
    Register_inst193 = 32'h0;	// <stdin>:5909:17, :6103:7
    Register_inst194 = 32'h0;	// <stdin>:5909:17, :6104:7
    Register_inst195 = 32'h0;	// <stdin>:5909:17, :6105:7
    Register_inst196 = 32'h0;	// <stdin>:5909:17, :6106:7
    Register_inst197 = 32'h0;	// <stdin>:5909:17, :6107:7
    Register_inst198 = 32'h0;	// <stdin>:5909:17, :6108:7
    Register_inst199 = 32'h0;	// <stdin>:5909:17, :6109:7
    Register_inst200 = 32'h0;	// <stdin>:5909:17, :6110:7
    Register_inst201 = 32'h0;	// <stdin>:5909:17, :6111:7
    Register_inst202 = 32'h0;	// <stdin>:5909:17, :6112:7
    Register_inst203 = 32'h0;	// <stdin>:5909:17, :6113:7
    Register_inst204 = 32'h0;	// <stdin>:5909:17, :6114:7
    Register_inst205 = 32'h0;	// <stdin>:5909:17, :6115:7
    Register_inst206 = 32'h0;	// <stdin>:5909:17, :6116:7
    Register_inst207 = 32'h0;	// <stdin>:5909:17, :6117:7
    Register_inst208 = 32'h0;	// <stdin>:5909:17, :6118:7
    Register_inst209 = 32'h0;	// <stdin>:5909:17, :6119:7
    Register_inst210 = 32'h0;	// <stdin>:5909:17, :6120:7
    Register_inst211 = 32'h0;	// <stdin>:5909:17, :6121:7
    Register_inst212 = 32'h0;	// <stdin>:5909:17, :6122:7
    Register_inst213 = 32'h0;	// <stdin>:5909:17, :6123:7
    Register_inst214 = 32'h0;	// <stdin>:5909:17, :6124:7
    Register_inst215 = 32'h0;	// <stdin>:5909:17, :6125:7
    Register_inst216 = 32'h0;	// <stdin>:5909:17, :6126:7
    Register_inst217 = 32'h0;	// <stdin>:5909:17, :6127:7
    Register_inst218 = 32'h0;	// <stdin>:5909:17, :6128:7
    Register_inst219 = 32'h0;	// <stdin>:5909:17, :6129:7
    Register_inst220 = 32'h0;	// <stdin>:5909:17, :6130:7
    Register_inst221 = 32'h0;	// <stdin>:5909:17, :6131:7
    Register_inst222 = 32'h0;	// <stdin>:5909:17, :6132:7
    Register_inst223 = 32'h0;	// <stdin>:5909:17, :6133:7
    Register_inst224 = 32'h0;	// <stdin>:5909:17, :6134:7
    Register_inst225 = 32'h0;	// <stdin>:5909:17, :6135:7
    Register_inst226 = 32'h0;	// <stdin>:5909:17, :6136:7
    Register_inst227 = 32'h0;	// <stdin>:5909:17, :6137:7
    Register_inst228 = 32'h0;	// <stdin>:5909:17, :6138:7
    Register_inst229 = 32'h0;	// <stdin>:5909:17, :6139:7
    Register_inst230 = 32'h0;	// <stdin>:5909:17, :6140:7
    Register_inst231 = 32'h0;	// <stdin>:5909:17, :6141:7
    Register_inst232 = 32'h0;	// <stdin>:5909:17, :6142:7
    Register_inst233 = 32'h0;	// <stdin>:5909:17, :6143:7
    Register_inst234 = 32'h0;	// <stdin>:5909:17, :6144:7
    Register_inst235 = 32'h0;	// <stdin>:5909:17, :6145:7
    Register_inst236 = 32'h0;	// <stdin>:5909:17, :6146:7
    Register_inst237 = 32'h0;	// <stdin>:5909:17, :6147:7
    Register_inst238 = 32'h0;	// <stdin>:5909:17, :6148:7
    Register_inst239 = 32'h0;	// <stdin>:5909:17, :6149:7
    Register_inst240 = 32'h0;	// <stdin>:5909:17, :6150:7
    Register_inst241 = 32'h0;	// <stdin>:5909:17, :6151:7
    Register_inst242 = 32'h0;	// <stdin>:5909:17, :6152:7
    Register_inst243 = 32'h0;	// <stdin>:5909:17, :6153:7
    Register_inst244 = 32'h0;	// <stdin>:5909:17, :6154:7
    Register_inst245 = 32'h0;	// <stdin>:5909:17, :6155:7
    Register_inst246 = 32'h0;	// <stdin>:5909:17, :6156:7
    Register_inst247 = 32'h0;	// <stdin>:5909:17, :6157:7
    Register_inst248 = 32'h0;	// <stdin>:5909:17, :6158:7
    Register_inst249 = 32'h0;	// <stdin>:5909:17, :6159:7
    Register_inst250 = 32'h0;	// <stdin>:5909:17, :6160:7
    Register_inst251 = 32'h0;	// <stdin>:5909:17, :6161:7
    Register_inst252 = 32'h0;	// <stdin>:5909:17, :6162:7
    Register_inst253 = 32'h0;	// <stdin>:5909:17, :6163:7
    Register_inst254 = 32'h0;	// <stdin>:5909:17, :6164:7
    Register_inst255 = 32'h0;	// <stdin>:5909:17, :6165:7
  end // initial
  assign _T = Register_inst255;	// <stdin>:6167:13
  wire [255:0][31:0] _tmp = {{_T_254}, {_T_253}, {_T_252}, {_T_251}, {_T_250}, {_T_249}, {_T_248}, {_T_247}, {_T_246}, {_T_245}, {_T_244}, {_T_243}, {_T_242}, {_T_241}, {_T_240}, {_T_239}, {_T_238}, {_T_237}, {_T_236}, {_T_235}, {_T_234}, {_T_233}, {_T_232}, {_T_231}, {_T_230}, {_T_229}, {_T_228}, {_T_227}, {_T_226}, {_T_225}, {_T_224}, {_T_223}, {_T_222}, {_T_221}, {_T_220}, {_T_219}, {_T_218}, {_T_217}, {_T_216}, {_T_215}, {_T_214}, {_T_213}, {_T_212}, {_T_211}, {_T_210}, {_T_209}, {_T_208}, {_T_207}, {_T_206}, {_T_205}, {_T_204}, {_T_203}, {_T_202}, {_T_201}, {_T_200}, {_T_199}, {_T_198}, {_T_197}, {_T_196}, {_T_195}, {_T_194}, {_T_193}, {_T_192}, {_T_191}, {_T_190}, {_T_189}, {_T_188}, {_T_187}, {_T_186}, {_T_185}, {_T_184}, {_T_183}, {_T_182}, {_T_181}, {_T_180}, {_T_179}, {_T_178}, {_T_177}, {_T_176}, {_T_175}, {_T_174}, {_T_173}, {_T_172}, {_T_171}, {_T_170}, {_T_169}, {_T_168}, {_T_167}, {_T_166}, {_T_165}, {_T_164}, {_T_163}, {_T_162}, {_T_161}, {_T_160}, {_T_159}, {_T_158}, {_T_157}, {_T_156}, {_T_155}, {_T_154}, {_T_153}, {_T_152}, {_T_151}, {_T_150}, {_T_149}, {_T_148}, {_T_147}, {_T_146}, {_T_145}, {_T_144}, {_T_143}, {_T_142}, {_T_141}, {_T_140}, {_T_139}, {_T_138}, {_T_137}, {_T_136}, {_T_135}, {_T_134}, {_T_133}, {_T_132}, {_T_131}, {_T_130}, {_T_129}, {_T_128}, {_T_127}, {_T_126}, {_T_125}, {_T_124}, {_T_123}, {_T_122}, {_T_121}, {_T_120}, {_T_119}, {_T_118}, {_T_117}, {_T_116}, {_T_115}, {_T_114}, {_T_113}, {_T_112}, {_T_111}, {_T_110}, {_T_109}, {_T_108}, {_T_107}, {_T_106}, {_T_105}, {_T_104}, {_T_103}, {_T_102}, {_T_101}, {_T_100}, {_T_99}, {_T_98}, {_T_97}, {_T_96}, {_T_95}, {_T_94}, {_T_93}, {_T_92}, {_T_91}, {_T_90}, {_T_89}, {_T_88}, {_T_87}, {_T_86}, {_T_85}, {_T_84}, {_T_83}, {_T_82}, {_T_81}, {_T_80}, {_T_79}, {_T_78}, {_T_77}, {_T_76}, {_T_75}, {_T_74}, {_T_73}, {_T_72}, {_T_71}, {_T_70}, {_T_69}, {_T_68}, {_T_67}, {_T_66}, {_T_65}, {_T_64}, {_T_63}, {_T_62}, {_T_61}, {_T_60}, {_T_59}, {_T_58}, {_T_57}, {_T_56}, {_T_55}, {_T_54}, {_T_53}, {_T_52}, {_T_51}, {_T_50}, {_T_49}, {_T_48}, {_T_47}, {_T_46}, {_T_45}, {_T_44}, {_T_43}, {_T_42}, {_T_41}, {_T_40}, {_T_39}, {_T_38}, {_T_37}, {_T_36}, {_T_35}, {_T_34}, {_T_33}, {_T_32}, {_T_31}, {_T_30}, {_T_29}, {_T_28}, {_T_27}, {_T_26}, {_T_25}, {_T_24}, {_T_23}, {_T_22}, {_T_21}, {_T_20}, {_T_19}, {_T_18}, {_T_17}, {_T_16}, {_T_15}, {_T_14}, {_T_13}, {_T_12}, {_T_11}, {_T_10}, {_T_9}, {_T_8}, {_T_7}, {_T_6}, {_T_5}, {_T_4}, {_T_3}, {_T_2}, {_T_1}, {_T_0}, {_T}};	// <stdin>:3352:10, :3360:11, :3368:11, :3376:11, :3384:11, :3392:11, :3400:11, :3408:11, :3416:11, :3424:11, :3432:11, :3440:11, :3448:11, :3456:11, :3464:12, :3472:12, :3480:12, :3488:12, :3496:12, :3504:12, :3512:12, :3520:12, :3528:12, :3536:12, :3544:12, :3552:12, :3560:12, :3568:12, :3576:12, :3584:12, :3592:12, :3600:12, :3608:12, :3616:12, :3624:12, :3632:12, :3640:12, :3648:12, :3656:12, :3664:12, :3672:12, :3680:12, :3688:12, :3696:12, :3704:12, :3712:12, :3720:12, :3728:12, :3736:12, :3744:12, :3752:12, :3760:12, :3768:12, :3776:12, :3784:12, :3792:12, :3800:12, :3808:12, :3816:12, :3824:12, :3832:12, :3840:12, :3848:12, :3856:12, :3864:12, :3872:12, :3880:12, :3888:12, :3896:12, :3904:12, :3912:12, :3920:12, :3928:12, :3936:12, :3944:12, :3952:12, :3960:12, :3968:12, :3976:12, :3984:12, :3992:12, :4000:12, :4008:12, :4016:12, :4024:12, :4032:12, :4040:12, :4048:12, :4056:12, :4064:12, :4072:12, :4080:12, :4088:12, :4096:12, :4104:12, :4112:12, :4120:12, :4128:12, :4136:12, :4144:12, :4152:12, :4160:12, :4168:12, :4176:12, :4184:12, :4192:12, :4200:12, :4208:12, :4216:12, :4224:12, :4232:12, :4240:12, :4248:12, :4256:12, :4264:12, :4272:12, :4280:12, :4288:12, :4296:12, :4304:12, :4312:12, :4320:12, :4328:12, :4336:12, :4344:12, :4352:12, :4360:12, :4368:12, :4376:12, :4384:12, :4392:12, :4400:12, :4408:12, :4416:12, :4424:12, :4432:12, :4440:12, :4448:12, :4456:12, :4464:12, :4472:12, :4480:12, :4488:13, :4496:13, :4504:13, :4512:13, :4520:13, :4528:13, :4536:13, :4544:13, :4552:13, :4560:13, :4568:13, :4576:13, :4584:13, :4592:13, :4600:13, :4608:13, :4616:13, :4624:13, :4632:13, :4640:13, :4648:13, :4656:13, :4664:13, :4672:13, :4680:13, :4688:13, :4696:13, :4704:13, :4712:13, :4720:13, :4728:13, :4736:13, :4744:13, :4752:13, :4760:13, :4768:13, :4776:13, :4784:13, :4792:13, :4800:13, :4808:13, :4816:13, :4824:13, :4832:13, :4840:13, :4848:13, :4856:13, :4864:13, :4872:13, :4880:13, :4888:13, :4896:13, :4904:13, :4912:13, :4920:13, :4928:13, :4936:13, :4944:13, :4952:13, :4960:13, :4968:13, :4976:13, :4984:13, :4992:13, :5000:13, :5008:13, :5016:13, :5024:13, :5032:13, :5040:13, :5048:13, :5056:13, :5064:13, :5072:13, :5080:13, :5088:13, :5096:13, :5104:13, :5112:13, :5120:13, :5128:13, :5136:13, :5144:13, :5152:13, :5160:13, :5168:13, :5176:13, :5184:13, :5192:13, :5200:13, :5208:13, :5216:13, :5224:13, :5232:13, :5240:13, :5248:13, :5256:13, :5264:13, :5272:13, :5280:13, :5288:13, :5296:13, :5304:13, :5312:13, :5320:13, :5328:13, :5336:13, :5344:13, :5352:13, :5360:13, :5368:13, :5376:13, :5384:13, :6167:13, :6168:13
  assign code_read_0_data = _tmp[code_read_0_addr];	// <stdin>:3352:10, :3360:11, :3368:11, :3376:11, :3384:11, :3392:11, :3400:11, :3408:11, :3416:11, :3424:11, :3432:11, :3440:11, :3448:11, :3456:11, :3464:12, :3472:12, :3480:12, :3488:12, :3496:12, :3504:12, :3512:12, :3520:12, :3528:12, :3536:12, :3544:12, :3552:12, :3560:12, :3568:12, :3576:12, :3584:12, :3592:12, :3600:12, :3608:12, :3616:12, :3624:12, :3632:12, :3640:12, :3648:12, :3656:12, :3664:12, :3672:12, :3680:12, :3688:12, :3696:12, :3704:12, :3712:12, :3720:12, :3728:12, :3736:12, :3744:12, :3752:12, :3760:12, :3768:12, :3776:12, :3784:12, :3792:12, :3800:12, :3808:12, :3816:12, :3824:12, :3832:12, :3840:12, :3848:12, :3856:12, :3864:12, :3872:12, :3880:12, :3888:12, :3896:12, :3904:12, :3912:12, :3920:12, :3928:12, :3936:12, :3944:12, :3952:12, :3960:12, :3968:12, :3976:12, :3984:12, :3992:12, :4000:12, :4008:12, :4016:12, :4024:12, :4032:12, :4040:12, :4048:12, :4056:12, :4064:12, :4072:12, :4080:12, :4088:12, :4096:12, :4104:12, :4112:12, :4120:12, :4128:12, :4136:12, :4144:12, :4152:12, :4160:12, :4168:12, :4176:12, :4184:12, :4192:12, :4200:12, :4208:12, :4216:12, :4224:12, :4232:12, :4240:12, :4248:12, :4256:12, :4264:12, :4272:12, :4280:12, :4288:12, :4296:12, :4304:12, :4312:12, :4320:12, :4328:12, :4336:12, :4344:12, :4352:12, :4360:12, :4368:12, :4376:12, :4384:12, :4392:12, :4400:12, :4408:12, :4416:12, :4424:12, :4432:12, :4440:12, :4448:12, :4456:12, :4464:12, :4472:12, :4480:12, :4488:13, :4496:13, :4504:13, :4512:13, :4520:13, :4528:13, :4536:13, :4544:13, :4552:13, :4560:13, :4568:13, :4576:13, :4584:13, :4592:13, :4600:13, :4608:13, :4616:13, :4624:13, :4632:13, :4640:13, :4648:13, :4656:13, :4664:13, :4672:13, :4680:13, :4688:13, :4696:13, :4704:13, :4712:13, :4720:13, :4728:13, :4736:13, :4744:13, :4752:13, :4760:13, :4768:13, :4776:13, :4784:13, :4792:13, :4800:13, :4808:13, :4816:13, :4824:13, :4832:13, :4840:13, :4848:13, :4856:13, :4864:13, :4872:13, :4880:13, :4888:13, :4896:13, :4904:13, :4912:13, :4920:13, :4928:13, :4936:13, :4944:13, :4952:13, :4960:13, :4968:13, :4976:13, :4984:13, :4992:13, :5000:13, :5008:13, :5016:13, :5024:13, :5032:13, :5040:13, :5048:13, :5056:13, :5064:13, :5072:13, :5080:13, :5088:13, :5096:13, :5104:13, :5112:13, :5120:13, :5128:13, :5136:13, :5144:13, :5152:13, :5160:13, :5168:13, :5176:13, :5184:13, :5192:13, :5200:13, :5208:13, :5216:13, :5224:13, :5232:13, :5240:13, :5248:13, :5256:13, :5264:13, :5272:13, :5280:13, :5288:13, :5296:13, :5304:13, :5312:13, :5320:13, :5328:13, :5336:13, :5344:13, :5352:13, :5360:13, :5368:13, :5376:13, :5384:13, :6167:13, :6169:13, :6170:5
endmodule

module Risc(
  input         is_write,
  input  [7:0]  write_addr,
  input  [31:0] write_data,
  input         boot, CLK, ASYNCRESET,
  output        valid,
  output [31:0] out);

  wire [31:0] _T;	// <stdin>:6238:11
  wire [7:0]  _T_0;	// <stdin>:6194:10
  wire [31:0] file_file_read_0_data;	// <stdin>:6221:54
  wire [31:0] file_file_read_1_data;	// <stdin>:6221:54
  wire [31:0] code_code_read_0_data;	// <stdin>:6196:30
  reg  [7:0]  Register_inst0;	// <stdin>:6186:23

  wire [7:0] _T_1 = ({{({{_T_0 + 8'h1}, {8'h0}})[boot]}, {_T_0}})[is_write];	// <stdin>:6177:14, :6178:14, :6181:10, :6182:10, :6183:10, :6184:10, :6185:10, :6194:10
  always @(posedge CLK)	// <stdin>:6187:5
    Register_inst0 <= _T_1;	// <stdin>:6188:7
  initial	// <stdin>:6190:5
    Register_inst0 = 8'h0;	// <stdin>:6191:18, :6192:7
  assign _T_0 = Register_inst0;	// <stdin>:6194:10
  wire struct packed {logic [31:0] data; logic [7:0] addr; } _T_2 = '{data: write_data, addr: write_addr};	// <stdin>:6195:10
  code code (	// <stdin>:6196:30
    .CLK              (CLK),
    .ASYNCRESET       (ASYNCRESET),
    .code_read_0_addr (_T_0),	// <stdin>:6194:10
    .write_0          (_T_2),
    .write_0_en       (is_write),
    .code_read_0_data (code_code_read_0_data)
  );
  wire [31:0] _T_3 = code_code_read_0_data;	// <stdin>:6196:30
  wire [31:0] _T_4 = code_code_read_0_data;	// <stdin>:6196:30
  wire [31:0] _T_5 = code_code_read_0_data;	// <stdin>:6196:30
  wire [31:0] _T_6 = code_code_read_0_data;	// <stdin>:6196:30
  wire [31:0] _T_7 = code_code_read_0_data;	// <stdin>:6196:30
  wire [31:0] _T_8 = code_code_read_0_data;	// <stdin>:6196:30
  wire [31:0] _T_9 = code_code_read_0_data;	// <stdin>:6196:30
  wire struct packed {logic [31:0] data; logic [7:0] addr; } _T_10 = '{data: _T, addr: (_T_9[23:16])};	// <stdin>:6216:11, :6217:11, :6238:11
  wire [31:0] _T_11 = code_code_read_0_data;	// <stdin>:6196:30
  file file (	// <stdin>:6221:54
    .CLK              (CLK),
    .ASYNCRESET       (ASYNCRESET),
    .file_read_0_addr (_T_7[15:8]),	// <stdin>:6214:11
    .file_read_1_addr (_T_8[7:0]),	// <stdin>:6215:11
    .write_0          (_T_10),
    .write_0_en       (~(&(_T_11[23:16]))),	// <stdin>:6218:11, :6219:11, :6220:11
    .file_read_0_data (file_file_read_0_data),
    .file_read_1_data (file_file_read_1_data)
  );
  wire [31:0] _T_12 = code_code_read_0_data;	// <stdin>:6196:30
  wire [31:0] _T_13 = code_code_read_0_data;	// <stdin>:6196:30
  wire [31:0] _T_14 = code_code_read_0_data;	// <stdin>:6196:30
  wire [31:0] _tmp = ({{32'h0}, {{24'h0, _T_4[15:8] << 8'h8 | _T_5[7:0]}}})[_T_6[31:24] == 8'h1];	// <stdin>:6173:15, :6174:14, :6175:15, :6178:14, :6205:11, :6206:11, :6207:11, :6208:11, :6209:11, :6210:11, :6211:11, :6212:11, :6213:11
  wire [31:0] _tmp_15 = ({{file_file_read_0_data}, {32'h0}})[_T_12[15:8] == 8'h0];	// <stdin>:6175:15, :6177:14, :6221:54, :6222:11, :6223:11, :6224:11, :6225:11
  wire [31:0] _tmp_16 = ({{file_file_read_1_data}, {32'h0}})[_T_13[7:0] == 8'h0];	// <stdin>:6175:15, :6177:14, :6221:54, :6226:11, :6227:11, :6228:11, :6229:11
  wire [31:0] _tmp_17 = ({{_tmp}, {_tmp_15 + _tmp_16}})[_T_14[31:24] == 8'h0];	// <stdin>:6177:14, :6230:11, :6231:11, :6232:11, :6233:11, :6234:11
  assign _T = ({{({{_tmp_17}, {32'h0}})[boot]}, {32'h0}})[is_write];	// <stdin>:6173:15, :6174:14, :6175:15, :6177:14, :6178:14, :6205:11, :6206:11, :6207:11, :6208:11, :6209:11, :6210:11, :6211:11, :6212:11, :6221:54, :6222:11, :6223:11, :6224:11, :6226:11, :6227:11, :6228:11, :6230:11, :6231:11, :6232:11, :6233:11, :6235:11, :6236:11, :6237:11, :6238:11
  wire _tmp_18 = ({{({{1'h0}, {1'h1}})[&(_T_3[23:16])]}, {1'h0}})[boot];	// <stdin>:6179:13, :6180:14, :6197:10, :6198:10, :6199:10, :6200:11, :6201:11, :6202:11
  assign valid = ({{_tmp_18}, {1'h0}})[is_write];	// <stdin>:6179:13, :6180:14, :6197:10, :6198:10, :6199:10, :6200:11, :6201:11, :6203:11, :6204:11, :6239:5
  assign out = _T;	// <stdin>:6238:11, :6239:5
endmodule

