module BasicALU(
  input  [3:0] a, b, opcode,
  output [3:0] out);

  wire [3:0] _tmp = ({{{3'h0, a == b}}, {{3'h0, a < b}}})[opcode == 4'h8];	// <stdin>:11:15, :12:14, :13:10, :14:10, :15:10, :16:10, :17:10, :18:10, :19:10
  wire [3:0] _tmp_0 = ({{({{_tmp}, {a - b}})[opcode == 4'h7]}, {a + b}})[opcode == 4'h6];	// <stdin>:9:14, :10:14, :20:10, :21:10, :22:10, :23:11, :24:11, :25:11, :26:11, :27:11
  wire [3:0] _tmp_1 = ({{({{_tmp_0}, {a - 4'h4}})[opcode == 4'h5]}, {a + 4'h4}})[opcode == 4'h4];	// <stdin>:7:14, :8:14, :28:16, :29:11, :30:11, :31:11, :32:11, :33:11, :34:11, :35:11, :36:11
  wire [3:0] _tmp_2 = ({{({{_tmp_1}, {a - 4'h1}})[opcode == 4'h3]}, {a + 4'h1}})[opcode == 4'h2];	// <stdin>:4:14, :5:14, :6:14, :37:16, :38:11, :39:11, :40:11, :41:11, :42:11, :43:11, :44:11, :45:11
  assign out = ({{({{_tmp_2}, {b}})[opcode == 4'h1]}, {a}})[opcode == 4'h0];	// <stdin>:3:14, :4:14, :5:14, :6:14, :7:14, :8:14, :9:14, :10:14, :11:15, :12:14, :13:10, :14:10, :15:10, :16:10, :17:10, :18:10, :20:10, :21:10, :22:10, :23:11, :24:11, :25:11, :26:11, :28:16, :29:11, :30:11, :31:11, :32:11, :33:11, :34:11, :35:11, :37:16, :38:11, :39:11, :40:11, :41:11, :42:11, :43:11, :44:11, :46:11, :47:11, :48:11, :49:11, :50:11, :51:11, :52:5
endmodule

