    module mod #(parameter KRATOS_INSTANCE_ID = 32'h0)
    (
        input I
    );

    endmodule   // mod
