module coreir_sgt #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output out
);
  assign out = $signed(in0) > $signed(in1);
endmodule

module TestBinary (
    input [6:0] I0,
    input [6:0] I1,
    output O
);
wire [6:0] magma_Bits_7_sgt_inst0_in0;
wire [6:0] magma_Bits_7_sgt_inst0_in1;
wire magma_Bits_7_sgt_inst0_out;
assign magma_Bits_7_sgt_inst0_in0 = I0;
assign magma_Bits_7_sgt_inst0_in1 = I1;
coreir_sgt #(
    .width(7)
) magma_Bits_7_sgt_inst0 (
    .in0(magma_Bits_7_sgt_inst0_in0),
    .in1(magma_Bits_7_sgt_inst0_in1),
    .out(magma_Bits_7_sgt_inst0_out)
);
assign O = magma_Bits_7_sgt_inst0_out;
endmodule

