module mantle_liftArrT__t_0Bit_1Bit21 (
    input in__0,
    input [1:0] in__1,
    output out_0__0,
    output [1:0] out_0__1
);
assign out_0__0 = in__0;
assign out_0__1 = in__1;
endmodule

module mantle_concatNArrT__Ns1__t_child_0BitIn_1BitIn2 (
    input in0_0__0,
    input [1:0] in0_0__1,
    output out_0__0,
    output [1:0] out_0__1
);
assign out_0__0 = in0_0__0;
assign out_0__1 = in0_0__1;
endmodule

module mantle_concatNArrT__Ns13__t_child_0BitIn_1BitIn2 (
    input in0_0__0,
    input [1:0] in0_0__1,
    input in1_0__0,
    input [1:0] in1_0__1,
    input in1_1__0,
    input [1:0] in1_1__1,
    input in1_2__0,
    input [1:0] in1_2__1,
    output out_0__0,
    output [1:0] out_0__1,
    output out_1__0,
    output [1:0] out_1__1,
    output out_2__0,
    output [1:0] out_2__1,
    output out_3__0,
    output [1:0] out_3__1
);
assign out_0__0 = in0_0__0;
assign out_0__1 = in0_0__1;
assign out_1__0 = in1_0__0;
assign out_1__1 = in1_0__1;
assign out_2__0 = in1_1__0;
assign out_2__1 = in1_1__1;
assign out_3__0 = in1_2__0;
assign out_3__1 = in1_2__1;
endmodule

module mantle_concatNArrT__Ns12__t_child_0BitIn_1BitIn2 (
    input in0_0__0,
    input [1:0] in0_0__1,
    input in1_0__0,
    input [1:0] in1_0__1,
    input in1_1__0,
    input [1:0] in1_1__1,
    output out_0__0,
    output [1:0] out_0__1,
    output out_1__0,
    output [1:0] out_1__1,
    output out_2__0,
    output [1:0] out_2__1
);
assign out_0__0 = in0_0__0;
assign out_0__1 = in0_0__1;
assign out_1__0 = in1_0__0;
assign out_1__1 = in1_0__1;
assign out_2__0 = in1_1__0;
assign out_2__1 = in1_1__1;
endmodule

module mantle_concatNArrT__Ns11__t_child_0BitIn_1BitIn2 (
    input in0_0__0,
    input [1:0] in0_0__1,
    input in1_0__0,
    input [1:0] in1_0__1,
    output out_0__0,
    output [1:0] out_0__1,
    output out_1__0,
    output [1:0] out_1__1
);
assign out_0__0 = in0_0__0;
assign out_0__1 = in0_0__1;
assign out_1__0 = in1_0__0;
assign out_1__1 = in1_0__1;
endmodule

module Foo (
    input I_0__0,
    input [1:0] I_0__1,
    input I_1__0,
    input [1:0] I_1__1,
    input I_2__0,
    input [1:0] I_2__1,
    input I_3__0,
    input [1:0] I_3__1,
    output O_0__0,
    output [1:0] O_0__1,
    output O_1__0,
    output [1:0] O_1__1,
    output O_2__0,
    output [1:0] O_2__1,
    output O_3__0,
    output [1:0] O_3__1
);
wire ConcatN_inst0_out_0__0;
wire [1:0] ConcatN_inst0_out_0__1;
wire ConcatN_inst0_out_1__0;
wire [1:0] ConcatN_inst0_out_1__1;
wire ConcatN_inst0_out_2__0;
wire [1:0] ConcatN_inst0_out_2__1;
wire ConcatN_inst0_out_3__0;
wire [1:0] ConcatN_inst0_out_3__1;
wire ConcatN_inst1_out_0__0;
wire [1:0] ConcatN_inst1_out_0__1;
wire ConcatN_inst1_out_1__0;
wire [1:0] ConcatN_inst1_out_1__1;
wire ConcatN_inst1_out_2__0;
wire [1:0] ConcatN_inst1_out_2__1;
wire ConcatN_inst2_out_0__0;
wire [1:0] ConcatN_inst2_out_0__1;
wire ConcatN_inst2_out_1__0;
wire [1:0] ConcatN_inst2_out_1__1;
wire ConcatN_inst3_out_0__0;
wire [1:0] ConcatN_inst3_out_0__1;
wire Lift_inst0_out_0__0;
wire [1:0] Lift_inst0_out_0__1;
wire Lift_inst1_out_0__0;
wire [1:0] Lift_inst1_out_0__1;
wire Lift_inst2_out_0__0;
wire [1:0] Lift_inst2_out_0__1;
wire Lift_inst3_out_0__0;
wire [1:0] Lift_inst3_out_0__1;
mantle_concatNArrT__Ns13__t_child_0BitIn_1BitIn2 ConcatN_inst0 (
    .in0_0__0(Lift_inst0_out_0__0),
    .in0_0__1(Lift_inst0_out_0__1),
    .in1_0__0(ConcatN_inst1_out_0__0),
    .in1_0__1(ConcatN_inst1_out_0__1),
    .in1_1__0(ConcatN_inst1_out_1__0),
    .in1_1__1(ConcatN_inst1_out_1__1),
    .in1_2__0(ConcatN_inst1_out_2__0),
    .in1_2__1(ConcatN_inst1_out_2__1),
    .out_0__0(ConcatN_inst0_out_0__0),
    .out_0__1(ConcatN_inst0_out_0__1),
    .out_1__0(ConcatN_inst0_out_1__0),
    .out_1__1(ConcatN_inst0_out_1__1),
    .out_2__0(ConcatN_inst0_out_2__0),
    .out_2__1(ConcatN_inst0_out_2__1),
    .out_3__0(ConcatN_inst0_out_3__0),
    .out_3__1(ConcatN_inst0_out_3__1)
);
mantle_concatNArrT__Ns12__t_child_0BitIn_1BitIn2 ConcatN_inst1 (
    .in0_0__0(Lift_inst1_out_0__0),
    .in0_0__1(Lift_inst1_out_0__1),
    .in1_0__0(ConcatN_inst2_out_0__0),
    .in1_0__1(ConcatN_inst2_out_0__1),
    .in1_1__0(ConcatN_inst2_out_1__0),
    .in1_1__1(ConcatN_inst2_out_1__1),
    .out_0__0(ConcatN_inst1_out_0__0),
    .out_0__1(ConcatN_inst1_out_0__1),
    .out_1__0(ConcatN_inst1_out_1__0),
    .out_1__1(ConcatN_inst1_out_1__1),
    .out_2__0(ConcatN_inst1_out_2__0),
    .out_2__1(ConcatN_inst1_out_2__1)
);
mantle_concatNArrT__Ns11__t_child_0BitIn_1BitIn2 ConcatN_inst2 (
    .in0_0__0(Lift_inst2_out_0__0),
    .in0_0__1(Lift_inst2_out_0__1),
    .in1_0__0(ConcatN_inst3_out_0__0),
    .in1_0__1(ConcatN_inst3_out_0__1),
    .out_0__0(ConcatN_inst2_out_0__0),
    .out_0__1(ConcatN_inst2_out_0__1),
    .out_1__0(ConcatN_inst2_out_1__0),
    .out_1__1(ConcatN_inst2_out_1__1)
);
mantle_concatNArrT__Ns1__t_child_0BitIn_1BitIn2 ConcatN_inst3 (
    .in0_0__0(Lift_inst3_out_0__0),
    .in0_0__1(Lift_inst3_out_0__1),
    .out_0__0(ConcatN_inst3_out_0__0),
    .out_0__1(ConcatN_inst3_out_0__1)
);
mantle_liftArrT__t_0Bit_1Bit21 Lift_inst0 (
    .in__0(I_3__0),
    .in__1(I_0__1),
    .out_0__0(Lift_inst0_out_0__0),
    .out_0__1(Lift_inst0_out_0__1)
);
mantle_liftArrT__t_0Bit_1Bit21 Lift_inst1 (
    .in__0(I_2__0),
    .in__1(I_1__1),
    .out_0__0(Lift_inst1_out_0__0),
    .out_0__1(Lift_inst1_out_0__1)
);
mantle_liftArrT__t_0Bit_1Bit21 Lift_inst2 (
    .in__0(I_1__0),
    .in__1(I_2__1),
    .out_0__0(Lift_inst2_out_0__0),
    .out_0__1(Lift_inst2_out_0__1)
);
mantle_liftArrT__t_0Bit_1Bit21 Lift_inst3 (
    .in__0(I_0__0),
    .in__1(I_3__1),
    .out_0__0(Lift_inst3_out_0__0),
    .out_0__1(Lift_inst3_out_0__1)
);
assign O_0__0 = ConcatN_inst0_out_0__0;
assign O_0__1 = ConcatN_inst0_out_0__1;
assign O_1__0 = ConcatN_inst0_out_1__0;
assign O_1__1 = ConcatN_inst0_out_1__1;
assign O_2__0 = ConcatN_inst0_out_2__0;
assign O_2__1 = ConcatN_inst0_out_2__1;
assign O_3__0 = ConcatN_inst0_out_3__0;
assign O_3__1 = ConcatN_inst0_out_3__1;
endmodule

