module mod5 #(parameter KRATOS_INSTANCE_ID = 17)
(
    input I
);

endmodule   // mod
