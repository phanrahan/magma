module simple_custom_verilog_name_custom_name(
  input  I,
  output O
);

  assign O = I;
endmodule

