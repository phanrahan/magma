module ByteSelector(
  input  [31:0] I,
  input  [1:0]  offset,
  output [7:0]  O);

  wire [7:0] _tmp = ({{({{I[31:24]}, {I[23:16]}})[offset == 2'h2]}, {I[15:8]}})[offset == 2'h1];	// <stdin>:4:14, :5:15, :6:10, :7:10, :8:10, :9:10, :10:10, :11:10, :12:10, :13:10, :14:10
  assign O = ({{_tmp}, {I[7:0]}})[offset == 2'h0];	// <stdin>:3:14, :4:14, :5:15, :6:10, :7:10, :8:10, :9:10, :10:10, :11:10, :12:10, :13:10, :15:10, :16:11, :17:11, :18:11, :19:5
endmodule

