module complex_aggregates_nested_array(
  input  [1:0][2:0][3:0] a,
  output [1:0][2:0][3:0] y);

  wire [3:0] _T = a[1'h0][2'h0];	// <stdin>:6:14, :7:14, :8:10, :9:10
  wire [3:0] _T_0 = a[1'h1][2'h2];	// <stdin>:4:15, :5:13, :11:10, :12:10
  wire [3:0] _T_1 = a[1'h0][2'h0];	// <stdin>:6:14, :7:14, :15:10, :16:10
  wire [3:0] _T_2 = a[1'h1][2'h2];	// <stdin>:4:15, :5:13, :18:11, :19:11
  wire [3:0] _T_3 = a[1'h0][2'h0];	// <stdin>:6:14, :7:14, :22:11, :23:11
  wire [3:0] _T_4 = a[1'h1][2'h2];	// <stdin>:4:15, :5:13, :25:11, :26:11
  wire [3:0] _T_5 = a[1'h0][2'h0];	// <stdin>:6:14, :7:14, :29:11, :30:11
  wire [3:0] _T_6 = a[1'h1][2'h2];	// <stdin>:4:15, :5:13, :32:11, :33:11
  wire [3:0] _T_7 = a[1'h0][2'h1];	// <stdin>:3:14, :7:14, :37:11, :38:11
  wire [3:0] _T_8 = a[1'h1][2'h1];	// <stdin>:3:14, :5:13, :40:11, :41:11
  wire [3:0] _T_9 = a[1'h0][2'h1];	// <stdin>:3:14, :7:14, :44:11, :45:11
  wire [3:0] _T_10 = a[1'h1][2'h1];	// <stdin>:3:14, :5:13, :47:11, :48:11
  wire [3:0] _T_11 = a[1'h0][2'h1];	// <stdin>:3:14, :7:14, :51:11, :52:11
  wire [3:0] _T_12 = a[1'h1][2'h1];	// <stdin>:3:14, :5:13, :54:11, :55:11
  wire [3:0] _T_13 = a[1'h0][2'h1];	// <stdin>:3:14, :7:14, :58:11, :59:11
  wire [3:0] _T_14 = a[1'h1][2'h1];	// <stdin>:3:14, :5:13, :61:11, :62:11
  wire [3:0] _T_15 = a[1'h0][2'h2];	// <stdin>:4:15, :7:14, :66:11, :67:11
  wire [3:0] _T_16 = a[1'h1][2'h0];	// <stdin>:5:13, :6:14, :69:11, :70:11
  wire [3:0] _T_17 = a[1'h0][2'h2];	// <stdin>:4:15, :7:14, :73:11, :74:11
  wire [3:0] _T_18 = a[1'h1][2'h0];	// <stdin>:5:13, :6:14, :76:11, :77:11
  wire [3:0] _T_19 = a[1'h0][2'h2];	// <stdin>:4:15, :7:14, :80:11, :81:11
  wire [3:0] _T_20 = a[1'h1][2'h0];	// <stdin>:5:13, :6:14, :83:11, :84:11
  wire [3:0] _T_21 = a[1'h0][2'h2];	// <stdin>:4:15, :7:14, :87:11, :88:11
  wire [3:0] _T_22 = a[1'h1][2'h0];	// <stdin>:5:13, :6:14, :90:11, :91:11
  wire [3:0] _T_23 = a[1'h1][2'h0];	// <stdin>:5:13, :6:14, :96:11, :97:11
  wire [3:0] _T_24 = a[1'h0][2'h2];	// <stdin>:4:15, :7:14, :99:11, :100:11
  wire [3:0] _T_25 = a[1'h1][2'h0];	// <stdin>:5:13, :6:14, :103:11, :104:11
  wire [3:0] _T_26 = a[1'h0][2'h2];	// <stdin>:4:15, :7:14, :106:11, :107:11
  wire [3:0] _T_27 = a[1'h1][2'h0];	// <stdin>:5:13, :6:14, :110:12, :111:12
  wire [3:0] _T_28 = a[1'h0][2'h2];	// <stdin>:4:15, :7:14, :113:12, :114:12
  wire [3:0] _T_29 = a[1'h1][2'h0];	// <stdin>:5:13, :6:14, :117:12, :118:12
  wire [3:0] _T_30 = a[1'h0][2'h2];	// <stdin>:4:15, :7:14, :120:12, :121:12
  wire [3:0] _T_31 = a[1'h1][2'h1];	// <stdin>:3:14, :5:13, :125:12, :126:12
  wire [3:0] _T_32 = a[1'h0][2'h1];	// <stdin>:3:14, :7:14, :128:12, :129:12
  wire [3:0] _T_33 = a[1'h1][2'h1];	// <stdin>:3:14, :5:13, :132:12, :133:12
  wire [3:0] _T_34 = a[1'h0][2'h1];	// <stdin>:3:14, :7:14, :135:12, :136:12
  wire [3:0] _T_35 = a[1'h1][2'h1];	// <stdin>:3:14, :5:13, :139:12, :140:12
  wire [3:0] _T_36 = a[1'h0][2'h1];	// <stdin>:3:14, :7:14, :142:12, :143:12
  wire [3:0] _T_37 = a[1'h1][2'h1];	// <stdin>:3:14, :5:13, :146:12, :147:12
  wire [3:0] _T_38 = a[1'h0][2'h1];	// <stdin>:3:14, :7:14, :149:12, :150:12
  wire [3:0] _T_39 = a[1'h1][2'h2];	// <stdin>:4:15, :5:13, :154:12, :155:12
  wire [3:0] _T_40 = a[1'h0][2'h0];	// <stdin>:6:14, :7:14, :157:12, :158:12
  wire [3:0] _T_41 = a[1'h1][2'h2];	// <stdin>:4:15, :5:13, :161:12, :162:12
  wire [3:0] _T_42 = a[1'h0][2'h0];	// <stdin>:6:14, :7:14, :164:12, :165:12
  wire [3:0] _T_43 = a[1'h1][2'h2];	// <stdin>:4:15, :5:13, :168:12, :169:12
  wire [3:0] _T_44 = a[1'h0][2'h0];	// <stdin>:6:14, :7:14, :171:12, :172:12
  wire [3:0] _T_45 = a[1'h1][2'h2];	// <stdin>:4:15, :5:13, :175:12, :176:12
  wire [3:0] _T_46 = a[1'h0][2'h0];	// <stdin>:6:14, :7:14, :178:12, :179:12
  wire [3:0] _tmp = {_T_45[3] | _T_46[0], _T_43[2] | _T_44[1], _T_41[1] | _T_42[2], _T_39[0] | _T_40[3]};	// <stdin>:156:12, :159:12, :160:12, :163:12, :166:12, :167:12, :170:12, :173:12, :174:12, :177:12, :180:12, :181:12, :182:12
  wire [3:0] _tmp_47 = {_T_37[3] | _T_38[0], _T_35[2] | _T_36[1], _T_33[1] | _T_34[2], _T_31[0] | _T_32[3]};	// <stdin>:127:12, :130:12, :131:12, :134:12, :137:12, :138:12, :141:12, :144:12, :145:12, :148:12, :151:12, :152:12, :153:12
  wire [3:0] _tmp_48 = {_T_29[3] | _T_30[0], _T_27[2] | _T_28[1], _T_25[1] | _T_26[2], _T_23[0] | _T_24[3]};	// <stdin>:98:11, :101:11, :102:11, :105:11, :108:12, :109:12, :112:12, :115:12, :116:12, :119:12, :122:12, :123:12, :124:12
  wire [3:0] _tmp_49 = {_T_21[3] | _T_22[0], _T_19[2] | _T_20[1], _T_17[1] | _T_18[2], _T_15[0] | _T_16[3]};	// <stdin>:68:11, :71:11, :72:11, :75:11, :78:11, :79:11, :82:11, :85:11, :86:11, :89:11, :92:11, :93:11, :94:11
  wire [3:0] _tmp_50 = {_T_13[3] | _T_14[0], _T_11[2] | _T_12[1], _T_9[1] | _T_10[2], _T_7[0] | _T_8[3]};	// <stdin>:39:11, :42:11, :43:11, :46:11, :49:11, :50:11, :53:11, :56:11, :57:11, :60:11, :63:11, :64:11, :65:11
  wire [3:0] _tmp_51 = {_T_5[3] | _T_6[0], _T_3[2] | _T_4[1], _T_1[1] | _T_2[2], _T[0] | _T_0[3]};	// <stdin>:10:10, :13:10, :14:10, :17:10, :20:11, :21:11, :24:11, :27:11, :28:11, :31:11, :34:11, :35:11, :36:11
  assign y = {{{{_tmp}, {_tmp_47}, {_tmp_48}}}, {{{_tmp_49}, {_tmp_50}, {_tmp_51}}}};	// <stdin>:10:10, :13:10, :14:10, :17:10, :20:11, :21:11, :24:11, :27:11, :28:11, :31:11, :34:11, :35:11, :39:11, :42:11, :43:11, :46:11, :49:11, :50:11, :53:11, :56:11, :57:11, :60:11, :63:11, :64:11, :68:11, :71:11, :72:11, :75:11, :78:11, :79:11, :82:11, :85:11, :86:11, :89:11, :92:11, :93:11, :95:11, :98:11, :101:11, :102:11, :105:11, :108:12, :109:12, :112:12, :115:12, :116:12, :119:12, :122:12, :123:12, :127:12, :130:12, :131:12, :134:12, :137:12, :138:12, :141:12, :144:12, :145:12, :148:12, :151:12, :152:12, :156:12, :159:12, :160:12, :163:12, :166:12, :167:12, :170:12, :173:12, :174:12, :177:12, :180:12, :181:12, :183:12, :184:12, :185:5
endmodule

