module mod2 #(parameter KRATOS_INSTANCE_ID = 24'd2)
(
    input I
);

endmodule   // mod
