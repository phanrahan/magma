module simple_smart_bits(
  input  [7:0] I,
  output [7:0] O
);

  assign O = I;
endmodule

