module TestCircuit (input [2:0] I_0_x, input [2:0] I_0_y, input [2:0] I_10_x, input [2:0] I_10_y, input [2:0] I_11_x, input [2:0] I_11_y, input [2:0] I_1_x, input [2:0] I_1_y, input [2:0] I_2_x, input [2:0] I_2_y, input [2:0] I_3_x, input [2:0] I_3_y, input [2:0] I_4_x, input [2:0] I_4_y, input [2:0] I_5_x, input [2:0] I_5_y, input [2:0] I_6_x, input [2:0] I_6_y, input [2:0] I_7_x, input [2:0] I_7_y, input [2:0] I_8_x, input [2:0] I_8_y, input [2:0] I_9_x, input [2:0] I_9_y, output [2:0] O_0_x, output [2:0] O_0_y, output [2:0] O_10_x, output [2:0] O_10_y, output [2:0] O_11_x, output [2:0] O_11_y, output [2:0] O_1_x, output [2:0] O_1_y, output [2:0] O_2_x, output [2:0] O_2_y, output [2:0] O_3_x, output [2:0] O_3_y, output [2:0] O_4_x, output [2:0] O_4_y, output [2:0] O_5_x, output [2:0] O_5_y, output [2:0] O_6_x, output [2:0] O_6_y, output [2:0] O_7_x, output [2:0] O_7_y, output [2:0] O_8_x, output [2:0] O_8_y, output [2:0] O_9_x, output [2:0] O_9_y);
assign O_0_x = I_0_x;
assign O_0_y = I_0_y;
assign O_10_x = I_10_x;
assign O_10_y = I_10_y;
assign O_11_x = I_11_x;
assign O_11_y = I_11_y;
assign O_1_x = I_1_x;
assign O_1_y = I_1_y;
assign O_2_x = I_2_x;
assign O_2_y = I_2_y;
assign O_3_x = I_3_x;
assign O_3_y = I_3_y;
assign O_4_x = I_4_x;
assign O_4_y = I_4_y;
assign O_5_x = I_5_x;
assign O_5_y = I_5_y;
assign O_6_x = I_6_x;
assign O_6_y = I_6_y;
assign O_7_x = I_7_x;
assign O_7_y = I_7_y;
assign O_8_x = I_8_x;
assign O_8_y = I_8_y;
assign O_9_x = I_9_x;
assign O_9_y = I_9_y;
endmodule

