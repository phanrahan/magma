module return_magma_tuple (input [1:0] I, output  O_0, output  O_1);
assign O_0 = I[0];
assign O_1 = I[1];
endmodule

