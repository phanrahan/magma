module basic_if (input [1:0] I_0, input  S_0, output  O);
assign O = I_0[1];
endmodule

