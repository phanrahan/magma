module top(a);
    input a;
endmodule
