module test_if_statement_basic (input [1:0] I, input  S, output  O);
assign O = I[0];
endmodule

