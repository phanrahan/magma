module return_py_tuple (input [1:0] I, output  O0, output  O1);
assign O0 = I[0];
assign O1 = I[1];
endmodule

