module file(	// <stdin>:1:1
  input                                                        CLK, ASYNCRESET,
  input  [7:0]                                                 file_read_0_addr,
  input  [7:0]                                                 file_read_1_addr,
  input  struct packed {logic [31:0] data; logic [7:0] addr; } write_0,
  input                                                        write_0_en,
  output [31:0]                                                file_read_0_data,
  output [31:0]                                                file_read_1_data);

  reg [31:0] Register_inst0;	// <stdin>:9:10
  reg [31:0] Register_inst1;	// <stdin>:25:11
  reg [31:0] Register_inst2;	// <stdin>:40:11
  reg [31:0] Register_inst3;	// <stdin>:55:11
  reg [31:0] Register_inst4;	// <stdin>:70:11
  reg [31:0] Register_inst5;	// <stdin>:85:11
  reg [31:0] Register_inst6;	// <stdin>:100:11
  reg [31:0] Register_inst7;	// <stdin>:115:11
  reg [31:0] Register_inst8;	// <stdin>:130:11
  reg [31:0] Register_inst9;	// <stdin>:145:11
  reg [31:0] Register_inst10;	// <stdin>:160:11
  reg [31:0] Register_inst11;	// <stdin>:175:11
  reg [31:0] Register_inst12;	// <stdin>:190:11
  reg [31:0] Register_inst13;	// <stdin>:205:12
  reg [31:0] Register_inst14;	// <stdin>:220:12
  reg [31:0] Register_inst15;	// <stdin>:235:12
  reg [31:0] Register_inst16;	// <stdin>:250:12
  reg [31:0] Register_inst17;	// <stdin>:265:12
  reg [31:0] Register_inst18;	// <stdin>:280:12
  reg [31:0] Register_inst19;	// <stdin>:295:12
  reg [31:0] Register_inst20;	// <stdin>:310:12
  reg [31:0] Register_inst21;	// <stdin>:325:12
  reg [31:0] Register_inst22;	// <stdin>:340:12
  reg [31:0] Register_inst23;	// <stdin>:355:12
  reg [31:0] Register_inst24;	// <stdin>:370:12
  reg [31:0] Register_inst25;	// <stdin>:385:12
  reg [31:0] Register_inst26;	// <stdin>:400:12
  reg [31:0] Register_inst27;	// <stdin>:415:12
  reg [31:0] Register_inst28;	// <stdin>:430:12
  reg [31:0] Register_inst29;	// <stdin>:445:12
  reg [31:0] Register_inst30;	// <stdin>:460:12
  reg [31:0] Register_inst31;	// <stdin>:475:12
  reg [31:0] Register_inst32;	// <stdin>:490:12
  reg [31:0] Register_inst33;	// <stdin>:505:12
  reg [31:0] Register_inst34;	// <stdin>:520:12
  reg [31:0] Register_inst35;	// <stdin>:535:12
  reg [31:0] Register_inst36;	// <stdin>:550:12
  reg [31:0] Register_inst37;	// <stdin>:565:12
  reg [31:0] Register_inst38;	// <stdin>:580:12
  reg [31:0] Register_inst39;	// <stdin>:595:12
  reg [31:0] Register_inst40;	// <stdin>:610:12
  reg [31:0] Register_inst41;	// <stdin>:625:12
  reg [31:0] Register_inst42;	// <stdin>:640:12
  reg [31:0] Register_inst43;	// <stdin>:655:12
  reg [31:0] Register_inst44;	// <stdin>:670:12
  reg [31:0] Register_inst45;	// <stdin>:685:12
  reg [31:0] Register_inst46;	// <stdin>:700:12
  reg [31:0] Register_inst47;	// <stdin>:715:12
  reg [31:0] Register_inst48;	// <stdin>:730:12
  reg [31:0] Register_inst49;	// <stdin>:745:12
  reg [31:0] Register_inst50;	// <stdin>:760:12
  reg [31:0] Register_inst51;	// <stdin>:775:12
  reg [31:0] Register_inst52;	// <stdin>:790:12
  reg [31:0] Register_inst53;	// <stdin>:805:12
  reg [31:0] Register_inst54;	// <stdin>:820:12
  reg [31:0] Register_inst55;	// <stdin>:835:12
  reg [31:0] Register_inst56;	// <stdin>:850:12
  reg [31:0] Register_inst57;	// <stdin>:865:12
  reg [31:0] Register_inst58;	// <stdin>:880:12
  reg [31:0] Register_inst59;	// <stdin>:895:12
  reg [31:0] Register_inst60;	// <stdin>:910:12
  reg [31:0] Register_inst61;	// <stdin>:925:12
  reg [31:0] Register_inst62;	// <stdin>:940:12
  reg [31:0] Register_inst63;	// <stdin>:955:12
  reg [31:0] Register_inst64;	// <stdin>:970:12
  reg [31:0] Register_inst65;	// <stdin>:985:12
  reg [31:0] Register_inst66;	// <stdin>:1000:12
  reg [31:0] Register_inst67;	// <stdin>:1015:12
  reg [31:0] Register_inst68;	// <stdin>:1030:12
  reg [31:0] Register_inst69;	// <stdin>:1045:12
  reg [31:0] Register_inst70;	// <stdin>:1060:12
  reg [31:0] Register_inst71;	// <stdin>:1075:12
  reg [31:0] Register_inst72;	// <stdin>:1090:12
  reg [31:0] Register_inst73;	// <stdin>:1105:12
  reg [31:0] Register_inst74;	// <stdin>:1120:12
  reg [31:0] Register_inst75;	// <stdin>:1135:12
  reg [31:0] Register_inst76;	// <stdin>:1150:12
  reg [31:0] Register_inst77;	// <stdin>:1165:12
  reg [31:0] Register_inst78;	// <stdin>:1180:12
  reg [31:0] Register_inst79;	// <stdin>:1195:12
  reg [31:0] Register_inst80;	// <stdin>:1210:12
  reg [31:0] Register_inst81;	// <stdin>:1225:12
  reg [31:0] Register_inst82;	// <stdin>:1240:12
  reg [31:0] Register_inst83;	// <stdin>:1255:12
  reg [31:0] Register_inst84;	// <stdin>:1270:12
  reg [31:0] Register_inst85;	// <stdin>:1285:12
  reg [31:0] Register_inst86;	// <stdin>:1300:12
  reg [31:0] Register_inst87;	// <stdin>:1315:12
  reg [31:0] Register_inst88;	// <stdin>:1330:12
  reg [31:0] Register_inst89;	// <stdin>:1345:12
  reg [31:0] Register_inst90;	// <stdin>:1360:12
  reg [31:0] Register_inst91;	// <stdin>:1375:12
  reg [31:0] Register_inst92;	// <stdin>:1390:12
  reg [31:0] Register_inst93;	// <stdin>:1405:12
  reg [31:0] Register_inst94;	// <stdin>:1420:12
  reg [31:0] Register_inst95;	// <stdin>:1435:12
  reg [31:0] Register_inst96;	// <stdin>:1450:12
  reg [31:0] Register_inst97;	// <stdin>:1465:12
  reg [31:0] Register_inst98;	// <stdin>:1480:12
  reg [31:0] Register_inst99;	// <stdin>:1495:12
  reg [31:0] Register_inst100;	// <stdin>:1510:12
  reg [31:0] Register_inst101;	// <stdin>:1525:12
  reg [31:0] Register_inst102;	// <stdin>:1540:12
  reg [31:0] Register_inst103;	// <stdin>:1555:12
  reg [31:0] Register_inst104;	// <stdin>:1570:12
  reg [31:0] Register_inst105;	// <stdin>:1585:12
  reg [31:0] Register_inst106;	// <stdin>:1600:12
  reg [31:0] Register_inst107;	// <stdin>:1615:12
  reg [31:0] Register_inst108;	// <stdin>:1630:12
  reg [31:0] Register_inst109;	// <stdin>:1645:12
  reg [31:0] Register_inst110;	// <stdin>:1660:12
  reg [31:0] Register_inst111;	// <stdin>:1675:12
  reg [31:0] Register_inst112;	// <stdin>:1690:12
  reg [31:0] Register_inst113;	// <stdin>:1705:12
  reg [31:0] Register_inst114;	// <stdin>:1720:12
  reg [31:0] Register_inst115;	// <stdin>:1735:12
  reg [31:0] Register_inst116;	// <stdin>:1750:12
  reg [31:0] Register_inst117;	// <stdin>:1765:12
  reg [31:0] Register_inst118;	// <stdin>:1780:12
  reg [31:0] Register_inst119;	// <stdin>:1795:12
  reg [31:0] Register_inst120;	// <stdin>:1810:12
  reg [31:0] Register_inst121;	// <stdin>:1825:12
  reg [31:0] Register_inst122;	// <stdin>:1840:12
  reg [31:0] Register_inst123;	// <stdin>:1855:12
  reg [31:0] Register_inst124;	// <stdin>:1870:12
  reg [31:0] Register_inst125;	// <stdin>:1885:12
  reg [31:0] Register_inst126;	// <stdin>:1900:12
  reg [31:0] Register_inst127;	// <stdin>:1915:12
  reg [31:0] Register_inst128;	// <stdin>:1930:12
  reg [31:0] Register_inst129;	// <stdin>:1945:12
  reg [31:0] Register_inst130;	// <stdin>:1960:12
  reg [31:0] Register_inst131;	// <stdin>:1975:12
  reg [31:0] Register_inst132;	// <stdin>:1990:12
  reg [31:0] Register_inst133;	// <stdin>:2005:12
  reg [31:0] Register_inst134;	// <stdin>:2020:12
  reg [31:0] Register_inst135;	// <stdin>:2035:12
  reg [31:0] Register_inst136;	// <stdin>:2050:12
  reg [31:0] Register_inst137;	// <stdin>:2065:12
  reg [31:0] Register_inst138;	// <stdin>:2080:12
  reg [31:0] Register_inst139;	// <stdin>:2095:12
  reg [31:0] Register_inst140;	// <stdin>:2110:12
  reg [31:0] Register_inst141;	// <stdin>:2125:12
  reg [31:0] Register_inst142;	// <stdin>:2140:13
  reg [31:0] Register_inst143;	// <stdin>:2155:13
  reg [31:0] Register_inst144;	// <stdin>:2170:13
  reg [31:0] Register_inst145;	// <stdin>:2185:13
  reg [31:0] Register_inst146;	// <stdin>:2200:13
  reg [31:0] Register_inst147;	// <stdin>:2215:13
  reg [31:0] Register_inst148;	// <stdin>:2230:13
  reg [31:0] Register_inst149;	// <stdin>:2245:13
  reg [31:0] Register_inst150;	// <stdin>:2260:13
  reg [31:0] Register_inst151;	// <stdin>:2275:13
  reg [31:0] Register_inst152;	// <stdin>:2290:13
  reg [31:0] Register_inst153;	// <stdin>:2305:13
  reg [31:0] Register_inst154;	// <stdin>:2320:13
  reg [31:0] Register_inst155;	// <stdin>:2335:13
  reg [31:0] Register_inst156;	// <stdin>:2350:13
  reg [31:0] Register_inst157;	// <stdin>:2365:13
  reg [31:0] Register_inst158;	// <stdin>:2380:13
  reg [31:0] Register_inst159;	// <stdin>:2395:13
  reg [31:0] Register_inst160;	// <stdin>:2410:13
  reg [31:0] Register_inst161;	// <stdin>:2425:13
  reg [31:0] Register_inst162;	// <stdin>:2440:13
  reg [31:0] Register_inst163;	// <stdin>:2455:13
  reg [31:0] Register_inst164;	// <stdin>:2470:13
  reg [31:0] Register_inst165;	// <stdin>:2485:13
  reg [31:0] Register_inst166;	// <stdin>:2500:13
  reg [31:0] Register_inst167;	// <stdin>:2515:13
  reg [31:0] Register_inst168;	// <stdin>:2530:13
  reg [31:0] Register_inst169;	// <stdin>:2545:13
  reg [31:0] Register_inst170;	// <stdin>:2560:13
  reg [31:0] Register_inst171;	// <stdin>:2575:13
  reg [31:0] Register_inst172;	// <stdin>:2590:13
  reg [31:0] Register_inst173;	// <stdin>:2605:13
  reg [31:0] Register_inst174;	// <stdin>:2620:13
  reg [31:0] Register_inst175;	// <stdin>:2635:13
  reg [31:0] Register_inst176;	// <stdin>:2650:13
  reg [31:0] Register_inst177;	// <stdin>:2665:13
  reg [31:0] Register_inst178;	// <stdin>:2680:13
  reg [31:0] Register_inst179;	// <stdin>:2695:13
  reg [31:0] Register_inst180;	// <stdin>:2710:13
  reg [31:0] Register_inst181;	// <stdin>:2725:13
  reg [31:0] Register_inst182;	// <stdin>:2740:13
  reg [31:0] Register_inst183;	// <stdin>:2755:13
  reg [31:0] Register_inst184;	// <stdin>:2770:13
  reg [31:0] Register_inst185;	// <stdin>:2785:13
  reg [31:0] Register_inst186;	// <stdin>:2800:13
  reg [31:0] Register_inst187;	// <stdin>:2815:13
  reg [31:0] Register_inst188;	// <stdin>:2830:13
  reg [31:0] Register_inst189;	// <stdin>:2845:13
  reg [31:0] Register_inst190;	// <stdin>:2860:13
  reg [31:0] Register_inst191;	// <stdin>:2875:13
  reg [31:0] Register_inst192;	// <stdin>:2890:13
  reg [31:0] Register_inst193;	// <stdin>:2905:13
  reg [31:0] Register_inst194;	// <stdin>:2920:13
  reg [31:0] Register_inst195;	// <stdin>:2935:13
  reg [31:0] Register_inst196;	// <stdin>:2950:13
  reg [31:0] Register_inst197;	// <stdin>:2965:13
  reg [31:0] Register_inst198;	// <stdin>:2980:13
  reg [31:0] Register_inst199;	// <stdin>:2995:13
  reg [31:0] Register_inst200;	// <stdin>:3010:13
  reg [31:0] Register_inst201;	// <stdin>:3025:13
  reg [31:0] Register_inst202;	// <stdin>:3040:13
  reg [31:0] Register_inst203;	// <stdin>:3055:13
  reg [31:0] Register_inst204;	// <stdin>:3070:13
  reg [31:0] Register_inst205;	// <stdin>:3085:13
  reg [31:0] Register_inst206;	// <stdin>:3100:13
  reg [31:0] Register_inst207;	// <stdin>:3115:13
  reg [31:0] Register_inst208;	// <stdin>:3130:13
  reg [31:0] Register_inst209;	// <stdin>:3145:13
  reg [31:0] Register_inst210;	// <stdin>:3160:13
  reg [31:0] Register_inst211;	// <stdin>:3175:13
  reg [31:0] Register_inst212;	// <stdin>:3190:13
  reg [31:0] Register_inst213;	// <stdin>:3205:13
  reg [31:0] Register_inst214;	// <stdin>:3220:13
  reg [31:0] Register_inst215;	// <stdin>:3235:13
  reg [31:0] Register_inst216;	// <stdin>:3250:13
  reg [31:0] Register_inst217;	// <stdin>:3265:13
  reg [31:0] Register_inst218;	// <stdin>:3280:13
  reg [31:0] Register_inst219;	// <stdin>:3295:13
  reg [31:0] Register_inst220;	// <stdin>:3310:13
  reg [31:0] Register_inst221;	// <stdin>:3325:13
  reg [31:0] Register_inst222;	// <stdin>:3340:13
  reg [31:0] Register_inst223;	// <stdin>:3355:13
  reg [31:0] Register_inst224;	// <stdin>:3370:13
  reg [31:0] Register_inst225;	// <stdin>:3385:13
  reg [31:0] Register_inst226;	// <stdin>:3400:13
  reg [31:0] Register_inst227;	// <stdin>:3415:13
  reg [31:0] Register_inst228;	// <stdin>:3430:13
  reg [31:0] Register_inst229;	// <stdin>:3445:13
  reg [31:0] Register_inst230;	// <stdin>:3460:13
  reg [31:0] Register_inst231;	// <stdin>:3475:13
  reg [31:0] Register_inst232;	// <stdin>:3490:13
  reg [31:0] Register_inst233;	// <stdin>:3505:13
  reg [31:0] Register_inst234;	// <stdin>:3520:13
  reg [31:0] Register_inst235;	// <stdin>:3535:13
  reg [31:0] Register_inst236;	// <stdin>:3550:13
  reg [31:0] Register_inst237;	// <stdin>:3565:13
  reg [31:0] Register_inst238;	// <stdin>:3580:13
  reg [31:0] Register_inst239;	// <stdin>:3595:13
  reg [31:0] Register_inst240;	// <stdin>:3610:13
  reg [31:0] Register_inst241;	// <stdin>:3625:13
  reg [31:0] Register_inst242;	// <stdin>:3640:13
  reg [31:0] Register_inst243;	// <stdin>:3655:13
  reg [31:0] Register_inst244;	// <stdin>:3670:13
  reg [31:0] Register_inst245;	// <stdin>:3685:13
  reg [31:0] Register_inst246;	// <stdin>:3700:13
  reg [31:0] Register_inst247;	// <stdin>:3715:13
  reg [31:0] Register_inst248;	// <stdin>:3730:13
  reg [31:0] Register_inst249;	// <stdin>:3745:13
  reg [31:0] Register_inst250;	// <stdin>:3760:13
  reg [31:0] Register_inst251;	// <stdin>:3775:13
  reg [31:0] Register_inst252;	// <stdin>:3790:13
  reg [31:0] Register_inst253;	// <stdin>:3805:13
  reg [31:0] Register_inst254;	// <stdin>:3820:13
  reg [31:0] Register_inst255;	// <stdin>:3835:13

  always_ff @(posedge CLK or posedge ASYNCRESET) begin	// <stdin>:3836:5
    if (ASYNCRESET) begin	// <stdin>:3836:5
      Register_inst0 <= 32'h0;	// <stdin>:13:9, :15:10
      Register_inst1 <= 32'h0;	// <stdin>:15:10, :29:9
      Register_inst2 <= 32'h0;	// <stdin>:15:10, :44:9
      Register_inst3 <= 32'h0;	// <stdin>:15:10, :59:9
      Register_inst4 <= 32'h0;	// <stdin>:15:10, :74:9
      Register_inst5 <= 32'h0;	// <stdin>:15:10, :89:9
      Register_inst6 <= 32'h0;	// <stdin>:15:10, :104:9
      Register_inst7 <= 32'h0;	// <stdin>:15:10, :119:9
      Register_inst8 <= 32'h0;	// <stdin>:15:10, :134:9
      Register_inst9 <= 32'h0;	// <stdin>:15:10, :149:9
      Register_inst10 <= 32'h0;	// <stdin>:15:10, :164:9
      Register_inst11 <= 32'h0;	// <stdin>:15:10, :179:9
      Register_inst12 <= 32'h0;	// <stdin>:15:10, :194:9
      Register_inst13 <= 32'h0;	// <stdin>:15:10, :209:9
      Register_inst14 <= 32'h0;	// <stdin>:15:10, :224:9
      Register_inst15 <= 32'h0;	// <stdin>:15:10, :239:9
      Register_inst16 <= 32'h0;	// <stdin>:15:10, :254:9
      Register_inst17 <= 32'h0;	// <stdin>:15:10, :269:9
      Register_inst18 <= 32'h0;	// <stdin>:15:10, :284:9
      Register_inst19 <= 32'h0;	// <stdin>:15:10, :299:9
      Register_inst20 <= 32'h0;	// <stdin>:15:10, :314:9
      Register_inst21 <= 32'h0;	// <stdin>:15:10, :329:9
      Register_inst22 <= 32'h0;	// <stdin>:15:10, :344:9
      Register_inst23 <= 32'h0;	// <stdin>:15:10, :359:9
      Register_inst24 <= 32'h0;	// <stdin>:15:10, :374:9
      Register_inst25 <= 32'h0;	// <stdin>:15:10, :389:9
      Register_inst26 <= 32'h0;	// <stdin>:15:10, :404:9
      Register_inst27 <= 32'h0;	// <stdin>:15:10, :419:9
      Register_inst28 <= 32'h0;	// <stdin>:15:10, :434:9
      Register_inst29 <= 32'h0;	// <stdin>:15:10, :449:9
      Register_inst30 <= 32'h0;	// <stdin>:15:10, :464:9
      Register_inst31 <= 32'h0;	// <stdin>:15:10, :479:9
      Register_inst32 <= 32'h0;	// <stdin>:15:10, :494:9
      Register_inst33 <= 32'h0;	// <stdin>:15:10, :509:9
      Register_inst34 <= 32'h0;	// <stdin>:15:10, :524:9
      Register_inst35 <= 32'h0;	// <stdin>:15:10, :539:9
      Register_inst36 <= 32'h0;	// <stdin>:15:10, :554:9
      Register_inst37 <= 32'h0;	// <stdin>:15:10, :569:9
      Register_inst38 <= 32'h0;	// <stdin>:15:10, :584:9
      Register_inst39 <= 32'h0;	// <stdin>:15:10, :599:9
      Register_inst40 <= 32'h0;	// <stdin>:15:10, :614:9
      Register_inst41 <= 32'h0;	// <stdin>:15:10, :629:9
      Register_inst42 <= 32'h0;	// <stdin>:15:10, :644:9
      Register_inst43 <= 32'h0;	// <stdin>:15:10, :659:9
      Register_inst44 <= 32'h0;	// <stdin>:15:10, :674:9
      Register_inst45 <= 32'h0;	// <stdin>:15:10, :689:9
      Register_inst46 <= 32'h0;	// <stdin>:15:10, :704:9
      Register_inst47 <= 32'h0;	// <stdin>:15:10, :719:9
      Register_inst48 <= 32'h0;	// <stdin>:15:10, :734:9
      Register_inst49 <= 32'h0;	// <stdin>:15:10, :749:9
      Register_inst50 <= 32'h0;	// <stdin>:15:10, :764:9
      Register_inst51 <= 32'h0;	// <stdin>:15:10, :779:9
      Register_inst52 <= 32'h0;	// <stdin>:15:10, :794:9
      Register_inst53 <= 32'h0;	// <stdin>:15:10, :809:9
      Register_inst54 <= 32'h0;	// <stdin>:15:10, :824:9
      Register_inst55 <= 32'h0;	// <stdin>:15:10, :839:9
      Register_inst56 <= 32'h0;	// <stdin>:15:10, :854:9
      Register_inst57 <= 32'h0;	// <stdin>:15:10, :869:9
      Register_inst58 <= 32'h0;	// <stdin>:15:10, :884:9
      Register_inst59 <= 32'h0;	// <stdin>:15:10, :899:9
      Register_inst60 <= 32'h0;	// <stdin>:15:10, :914:9
      Register_inst61 <= 32'h0;	// <stdin>:15:10, :929:9
      Register_inst62 <= 32'h0;	// <stdin>:15:10, :944:9
      Register_inst63 <= 32'h0;	// <stdin>:15:10, :959:9
      Register_inst64 <= 32'h0;	// <stdin>:15:10, :974:9
      Register_inst65 <= 32'h0;	// <stdin>:15:10, :989:9
      Register_inst66 <= 32'h0;	// <stdin>:15:10, :1004:9
      Register_inst67 <= 32'h0;	// <stdin>:15:10, :1019:9
      Register_inst68 <= 32'h0;	// <stdin>:15:10, :1034:9
      Register_inst69 <= 32'h0;	// <stdin>:15:10, :1049:9
      Register_inst70 <= 32'h0;	// <stdin>:15:10, :1064:9
      Register_inst71 <= 32'h0;	// <stdin>:15:10, :1079:9
      Register_inst72 <= 32'h0;	// <stdin>:15:10, :1094:9
      Register_inst73 <= 32'h0;	// <stdin>:15:10, :1109:9
      Register_inst74 <= 32'h0;	// <stdin>:15:10, :1124:9
      Register_inst75 <= 32'h0;	// <stdin>:15:10, :1139:9
      Register_inst76 <= 32'h0;	// <stdin>:15:10, :1154:9
      Register_inst77 <= 32'h0;	// <stdin>:15:10, :1169:9
      Register_inst78 <= 32'h0;	// <stdin>:15:10, :1184:9
      Register_inst79 <= 32'h0;	// <stdin>:15:10, :1199:9
      Register_inst80 <= 32'h0;	// <stdin>:15:10, :1214:9
      Register_inst81 <= 32'h0;	// <stdin>:15:10, :1229:9
      Register_inst82 <= 32'h0;	// <stdin>:15:10, :1244:9
      Register_inst83 <= 32'h0;	// <stdin>:15:10, :1259:9
      Register_inst84 <= 32'h0;	// <stdin>:15:10, :1274:9
      Register_inst85 <= 32'h0;	// <stdin>:15:10, :1289:9
      Register_inst86 <= 32'h0;	// <stdin>:15:10, :1304:9
      Register_inst87 <= 32'h0;	// <stdin>:15:10, :1319:9
      Register_inst88 <= 32'h0;	// <stdin>:15:10, :1334:9
      Register_inst89 <= 32'h0;	// <stdin>:15:10, :1349:9
      Register_inst90 <= 32'h0;	// <stdin>:15:10, :1364:9
      Register_inst91 <= 32'h0;	// <stdin>:15:10, :1379:9
      Register_inst92 <= 32'h0;	// <stdin>:15:10, :1394:9
      Register_inst93 <= 32'h0;	// <stdin>:15:10, :1409:9
      Register_inst94 <= 32'h0;	// <stdin>:15:10, :1424:9
      Register_inst95 <= 32'h0;	// <stdin>:15:10, :1439:9
      Register_inst96 <= 32'h0;	// <stdin>:15:10, :1454:9
      Register_inst97 <= 32'h0;	// <stdin>:15:10, :1469:9
      Register_inst98 <= 32'h0;	// <stdin>:15:10, :1484:9
      Register_inst99 <= 32'h0;	// <stdin>:15:10, :1499:9
      Register_inst100 <= 32'h0;	// <stdin>:15:10, :1514:9
      Register_inst101 <= 32'h0;	// <stdin>:15:10, :1529:9
      Register_inst102 <= 32'h0;	// <stdin>:15:10, :1544:9
      Register_inst103 <= 32'h0;	// <stdin>:15:10, :1559:9
      Register_inst104 <= 32'h0;	// <stdin>:15:10, :1574:9
      Register_inst105 <= 32'h0;	// <stdin>:15:10, :1589:9
      Register_inst106 <= 32'h0;	// <stdin>:15:10, :1604:9
      Register_inst107 <= 32'h0;	// <stdin>:15:10, :1619:9
      Register_inst108 <= 32'h0;	// <stdin>:15:10, :1634:9
      Register_inst109 <= 32'h0;	// <stdin>:15:10, :1649:9
      Register_inst110 <= 32'h0;	// <stdin>:15:10, :1664:9
      Register_inst111 <= 32'h0;	// <stdin>:15:10, :1679:9
      Register_inst112 <= 32'h0;	// <stdin>:15:10, :1694:9
      Register_inst113 <= 32'h0;	// <stdin>:15:10, :1709:9
      Register_inst114 <= 32'h0;	// <stdin>:15:10, :1724:9
      Register_inst115 <= 32'h0;	// <stdin>:15:10, :1739:9
      Register_inst116 <= 32'h0;	// <stdin>:15:10, :1754:9
      Register_inst117 <= 32'h0;	// <stdin>:15:10, :1769:9
      Register_inst118 <= 32'h0;	// <stdin>:15:10, :1784:9
      Register_inst119 <= 32'h0;	// <stdin>:15:10, :1799:9
      Register_inst120 <= 32'h0;	// <stdin>:15:10, :1814:9
      Register_inst121 <= 32'h0;	// <stdin>:15:10, :1829:9
      Register_inst122 <= 32'h0;	// <stdin>:15:10, :1844:9
      Register_inst123 <= 32'h0;	// <stdin>:15:10, :1859:9
      Register_inst124 <= 32'h0;	// <stdin>:15:10, :1874:9
      Register_inst125 <= 32'h0;	// <stdin>:15:10, :1889:9
      Register_inst126 <= 32'h0;	// <stdin>:15:10, :1904:9
      Register_inst127 <= 32'h0;	// <stdin>:15:10, :1919:9
      Register_inst128 <= 32'h0;	// <stdin>:15:10, :1934:9
      Register_inst129 <= 32'h0;	// <stdin>:15:10, :1949:9
      Register_inst130 <= 32'h0;	// <stdin>:15:10, :1964:9
      Register_inst131 <= 32'h0;	// <stdin>:15:10, :1979:9
      Register_inst132 <= 32'h0;	// <stdin>:15:10, :1994:9
      Register_inst133 <= 32'h0;	// <stdin>:15:10, :2009:9
      Register_inst134 <= 32'h0;	// <stdin>:15:10, :2024:9
      Register_inst135 <= 32'h0;	// <stdin>:15:10, :2039:9
      Register_inst136 <= 32'h0;	// <stdin>:15:10, :2054:9
      Register_inst137 <= 32'h0;	// <stdin>:15:10, :2069:9
      Register_inst138 <= 32'h0;	// <stdin>:15:10, :2084:9
      Register_inst139 <= 32'h0;	// <stdin>:15:10, :2099:9
      Register_inst140 <= 32'h0;	// <stdin>:15:10, :2114:9
      Register_inst141 <= 32'h0;	// <stdin>:15:10, :2129:9
      Register_inst142 <= 32'h0;	// <stdin>:15:10, :2144:9
      Register_inst143 <= 32'h0;	// <stdin>:15:10, :2159:9
      Register_inst144 <= 32'h0;	// <stdin>:15:10, :2174:9
      Register_inst145 <= 32'h0;	// <stdin>:15:10, :2189:9
      Register_inst146 <= 32'h0;	// <stdin>:15:10, :2204:9
      Register_inst147 <= 32'h0;	// <stdin>:15:10, :2219:9
      Register_inst148 <= 32'h0;	// <stdin>:15:10, :2234:9
      Register_inst149 <= 32'h0;	// <stdin>:15:10, :2249:9
      Register_inst150 <= 32'h0;	// <stdin>:15:10, :2264:9
      Register_inst151 <= 32'h0;	// <stdin>:15:10, :2279:9
      Register_inst152 <= 32'h0;	// <stdin>:15:10, :2294:9
      Register_inst153 <= 32'h0;	// <stdin>:15:10, :2309:9
      Register_inst154 <= 32'h0;	// <stdin>:15:10, :2324:9
      Register_inst155 <= 32'h0;	// <stdin>:15:10, :2339:9
      Register_inst156 <= 32'h0;	// <stdin>:15:10, :2354:9
      Register_inst157 <= 32'h0;	// <stdin>:15:10, :2369:9
      Register_inst158 <= 32'h0;	// <stdin>:15:10, :2384:9
      Register_inst159 <= 32'h0;	// <stdin>:15:10, :2399:9
      Register_inst160 <= 32'h0;	// <stdin>:15:10, :2414:9
      Register_inst161 <= 32'h0;	// <stdin>:15:10, :2429:9
      Register_inst162 <= 32'h0;	// <stdin>:15:10, :2444:9
      Register_inst163 <= 32'h0;	// <stdin>:15:10, :2459:9
      Register_inst164 <= 32'h0;	// <stdin>:15:10, :2474:9
      Register_inst165 <= 32'h0;	// <stdin>:15:10, :2489:9
      Register_inst166 <= 32'h0;	// <stdin>:15:10, :2504:9
      Register_inst167 <= 32'h0;	// <stdin>:15:10, :2519:9
      Register_inst168 <= 32'h0;	// <stdin>:15:10, :2534:9
      Register_inst169 <= 32'h0;	// <stdin>:15:10, :2549:9
      Register_inst170 <= 32'h0;	// <stdin>:15:10, :2564:9
      Register_inst171 <= 32'h0;	// <stdin>:15:10, :2579:9
      Register_inst172 <= 32'h0;	// <stdin>:15:10, :2594:9
      Register_inst173 <= 32'h0;	// <stdin>:15:10, :2609:9
      Register_inst174 <= 32'h0;	// <stdin>:15:10, :2624:9
      Register_inst175 <= 32'h0;	// <stdin>:15:10, :2639:9
      Register_inst176 <= 32'h0;	// <stdin>:15:10, :2654:9
      Register_inst177 <= 32'h0;	// <stdin>:15:10, :2669:9
      Register_inst178 <= 32'h0;	// <stdin>:15:10, :2684:9
      Register_inst179 <= 32'h0;	// <stdin>:15:10, :2699:9
      Register_inst180 <= 32'h0;	// <stdin>:15:10, :2714:9
      Register_inst181 <= 32'h0;	// <stdin>:15:10, :2729:9
      Register_inst182 <= 32'h0;	// <stdin>:15:10, :2744:9
      Register_inst183 <= 32'h0;	// <stdin>:15:10, :2759:9
      Register_inst184 <= 32'h0;	// <stdin>:15:10, :2774:9
      Register_inst185 <= 32'h0;	// <stdin>:15:10, :2789:9
      Register_inst186 <= 32'h0;	// <stdin>:15:10, :2804:9
      Register_inst187 <= 32'h0;	// <stdin>:15:10, :2819:9
      Register_inst188 <= 32'h0;	// <stdin>:15:10, :2834:9
      Register_inst189 <= 32'h0;	// <stdin>:15:10, :2849:9
      Register_inst190 <= 32'h0;	// <stdin>:15:10, :2864:9
      Register_inst191 <= 32'h0;	// <stdin>:15:10, :2879:9
      Register_inst192 <= 32'h0;	// <stdin>:15:10, :2894:9
      Register_inst193 <= 32'h0;	// <stdin>:15:10, :2909:9
      Register_inst194 <= 32'h0;	// <stdin>:15:10, :2924:9
      Register_inst195 <= 32'h0;	// <stdin>:15:10, :2939:9
      Register_inst196 <= 32'h0;	// <stdin>:15:10, :2954:9
      Register_inst197 <= 32'h0;	// <stdin>:15:10, :2969:9
      Register_inst198 <= 32'h0;	// <stdin>:15:10, :2984:9
      Register_inst199 <= 32'h0;	// <stdin>:15:10, :2999:9
      Register_inst200 <= 32'h0;	// <stdin>:15:10, :3014:9
      Register_inst201 <= 32'h0;	// <stdin>:15:10, :3029:9
      Register_inst202 <= 32'h0;	// <stdin>:15:10, :3044:9
      Register_inst203 <= 32'h0;	// <stdin>:15:10, :3059:9
      Register_inst204 <= 32'h0;	// <stdin>:15:10, :3074:9
      Register_inst205 <= 32'h0;	// <stdin>:15:10, :3089:9
      Register_inst206 <= 32'h0;	// <stdin>:15:10, :3104:9
      Register_inst207 <= 32'h0;	// <stdin>:15:10, :3119:9
      Register_inst208 <= 32'h0;	// <stdin>:15:10, :3134:9
      Register_inst209 <= 32'h0;	// <stdin>:15:10, :3149:9
      Register_inst210 <= 32'h0;	// <stdin>:15:10, :3164:9
      Register_inst211 <= 32'h0;	// <stdin>:15:10, :3179:9
      Register_inst212 <= 32'h0;	// <stdin>:15:10, :3194:9
      Register_inst213 <= 32'h0;	// <stdin>:15:10, :3209:9
      Register_inst214 <= 32'h0;	// <stdin>:15:10, :3224:9
      Register_inst215 <= 32'h0;	// <stdin>:15:10, :3239:9
      Register_inst216 <= 32'h0;	// <stdin>:15:10, :3254:9
      Register_inst217 <= 32'h0;	// <stdin>:15:10, :3269:9
      Register_inst218 <= 32'h0;	// <stdin>:15:10, :3284:9
      Register_inst219 <= 32'h0;	// <stdin>:15:10, :3299:9
      Register_inst220 <= 32'h0;	// <stdin>:15:10, :3314:9
      Register_inst221 <= 32'h0;	// <stdin>:15:10, :3329:9
      Register_inst222 <= 32'h0;	// <stdin>:15:10, :3344:9
      Register_inst223 <= 32'h0;	// <stdin>:15:10, :3359:9
      Register_inst224 <= 32'h0;	// <stdin>:15:10, :3374:9
      Register_inst225 <= 32'h0;	// <stdin>:15:10, :3389:9
      Register_inst226 <= 32'h0;	// <stdin>:15:10, :3404:9
      Register_inst227 <= 32'h0;	// <stdin>:15:10, :3419:9
      Register_inst228 <= 32'h0;	// <stdin>:15:10, :3434:9
      Register_inst229 <= 32'h0;	// <stdin>:15:10, :3449:9
      Register_inst230 <= 32'h0;	// <stdin>:15:10, :3464:9
      Register_inst231 <= 32'h0;	// <stdin>:15:10, :3479:9
      Register_inst232 <= 32'h0;	// <stdin>:15:10, :3494:9
      Register_inst233 <= 32'h0;	// <stdin>:15:10, :3509:9
      Register_inst234 <= 32'h0;	// <stdin>:15:10, :3524:9
      Register_inst235 <= 32'h0;	// <stdin>:15:10, :3539:9
      Register_inst236 <= 32'h0;	// <stdin>:15:10, :3554:9
      Register_inst237 <= 32'h0;	// <stdin>:15:10, :3569:9
      Register_inst238 <= 32'h0;	// <stdin>:15:10, :3584:9
      Register_inst239 <= 32'h0;	// <stdin>:15:10, :3599:9
      Register_inst240 <= 32'h0;	// <stdin>:15:10, :3614:9
      Register_inst241 <= 32'h0;	// <stdin>:15:10, :3629:9
      Register_inst242 <= 32'h0;	// <stdin>:15:10, :3644:9
      Register_inst243 <= 32'h0;	// <stdin>:15:10, :3659:9
      Register_inst244 <= 32'h0;	// <stdin>:15:10, :3674:9
      Register_inst245 <= 32'h0;	// <stdin>:15:10, :3689:9
      Register_inst246 <= 32'h0;	// <stdin>:15:10, :3704:9
      Register_inst247 <= 32'h0;	// <stdin>:15:10, :3719:9
      Register_inst248 <= 32'h0;	// <stdin>:15:10, :3734:9
      Register_inst249 <= 32'h0;	// <stdin>:15:10, :3749:9
      Register_inst250 <= 32'h0;	// <stdin>:15:10, :3764:9
      Register_inst251 <= 32'h0;	// <stdin>:15:10, :3779:9
      Register_inst252 <= 32'h0;	// <stdin>:15:10, :3794:9
      Register_inst253 <= 32'h0;	// <stdin>:15:10, :3809:9
      Register_inst254 <= 32'h0;	// <stdin>:15:10, :3824:9
      Register_inst255 <= 32'h0;	// <stdin>:15:10, :3839:9
    end
    else begin	// <stdin>:3836:5
      automatic logic [31:0]      _T_1 = write_0.data;	// <stdin>:2:10
      automatic logic [7:0]       _T_2 = write_0.addr;	// <stdin>:3:10
      automatic logic [1:0][31:0] _T_3 = {{Register_inst0}, {_T_1}};	// <stdin>:7:10, :19:10
      automatic logic [1:0][31:0] _T_4 = {{Register_inst1}, {_T_1}};	// <stdin>:23:11, :34:11
      automatic logic [1:0][31:0] _T_5 = {{Register_inst2}, {_T_1}};	// <stdin>:38:11, :49:11
      automatic logic [1:0][31:0] _T_6 = {{Register_inst3}, {_T_1}};	// <stdin>:53:11, :64:11
      automatic logic [1:0][31:0] _T_7 = {{Register_inst4}, {_T_1}};	// <stdin>:68:11, :79:11
      automatic logic [1:0][31:0] _T_8 = {{Register_inst5}, {_T_1}};	// <stdin>:83:11, :94:11
      automatic logic [1:0][31:0] _T_9 = {{Register_inst6}, {_T_1}};	// <stdin>:98:11, :109:11
      automatic logic [1:0][31:0] _T_10 = {{Register_inst7}, {_T_1}};	// <stdin>:113:11, :124:11
      automatic logic [1:0][31:0] _T_11 = {{Register_inst8}, {_T_1}};	// <stdin>:128:11, :139:11
      automatic logic [1:0][31:0] _T_12 = {{Register_inst9}, {_T_1}};	// <stdin>:143:11, :154:11
      automatic logic [1:0][31:0] _T_13 = {{Register_inst10}, {_T_1}};	// <stdin>:158:11, :169:11
      automatic logic [1:0][31:0] _T_14 = {{Register_inst11}, {_T_1}};	// <stdin>:173:11, :184:11
      automatic logic [1:0][31:0] _T_15 = {{Register_inst12}, {_T_1}};	// <stdin>:188:11, :199:11
      automatic logic [1:0][31:0] _T_16 = {{Register_inst13}, {_T_1}};	// <stdin>:203:11, :214:11
      automatic logic [1:0][31:0] _T_17 = {{Register_inst14}, {_T_1}};	// <stdin>:218:12, :229:12
      automatic logic [1:0][31:0] _T_18 = {{Register_inst15}, {_T_1}};	// <stdin>:233:12, :244:12
      automatic logic [1:0][31:0] _T_19 = {{Register_inst16}, {_T_1}};	// <stdin>:248:12, :259:12
      automatic logic [1:0][31:0] _T_20 = {{Register_inst17}, {_T_1}};	// <stdin>:263:12, :274:12
      automatic logic [1:0][31:0] _T_21 = {{Register_inst18}, {_T_1}};	// <stdin>:278:12, :289:12
      automatic logic [1:0][31:0] _T_22 = {{Register_inst19}, {_T_1}};	// <stdin>:293:12, :304:12
      automatic logic [1:0][31:0] _T_23 = {{Register_inst20}, {_T_1}};	// <stdin>:308:12, :319:12
      automatic logic [1:0][31:0] _T_24 = {{Register_inst21}, {_T_1}};	// <stdin>:323:12, :334:12
      automatic logic [1:0][31:0] _T_25 = {{Register_inst22}, {_T_1}};	// <stdin>:338:12, :349:12
      automatic logic [1:0][31:0] _T_26 = {{Register_inst23}, {_T_1}};	// <stdin>:353:12, :364:12
      automatic logic [1:0][31:0] _T_27 = {{Register_inst24}, {_T_1}};	// <stdin>:368:12, :379:12
      automatic logic [1:0][31:0] _T_28 = {{Register_inst25}, {_T_1}};	// <stdin>:383:12, :394:12
      automatic logic [1:0][31:0] _T_29 = {{Register_inst26}, {_T_1}};	// <stdin>:398:12, :409:12
      automatic logic [1:0][31:0] _T_30 = {{Register_inst27}, {_T_1}};	// <stdin>:413:12, :424:12
      automatic logic [1:0][31:0] _T_31 = {{Register_inst28}, {_T_1}};	// <stdin>:428:12, :439:12
      automatic logic [1:0][31:0] _T_32 = {{Register_inst29}, {_T_1}};	// <stdin>:443:12, :454:12
      automatic logic [1:0][31:0] _T_33 = {{Register_inst30}, {_T_1}};	// <stdin>:458:12, :469:12
      automatic logic [1:0][31:0] _T_34 = {{Register_inst31}, {_T_1}};	// <stdin>:473:12, :484:12
      automatic logic [1:0][31:0] _T_35 = {{Register_inst32}, {_T_1}};	// <stdin>:488:12, :499:12
      automatic logic [1:0][31:0] _T_36 = {{Register_inst33}, {_T_1}};	// <stdin>:503:12, :514:12
      automatic logic [1:0][31:0] _T_37 = {{Register_inst34}, {_T_1}};	// <stdin>:518:12, :529:12
      automatic logic [1:0][31:0] _T_38 = {{Register_inst35}, {_T_1}};	// <stdin>:533:12, :544:12
      automatic logic [1:0][31:0] _T_39 = {{Register_inst36}, {_T_1}};	// <stdin>:548:12, :559:12
      automatic logic [1:0][31:0] _T_40 = {{Register_inst37}, {_T_1}};	// <stdin>:563:12, :574:12
      automatic logic [1:0][31:0] _T_41 = {{Register_inst38}, {_T_1}};	// <stdin>:578:12, :589:12
      automatic logic [1:0][31:0] _T_42 = {{Register_inst39}, {_T_1}};	// <stdin>:593:12, :604:12
      automatic logic [1:0][31:0] _T_43 = {{Register_inst40}, {_T_1}};	// <stdin>:608:12, :619:12
      automatic logic [1:0][31:0] _T_44 = {{Register_inst41}, {_T_1}};	// <stdin>:623:12, :634:12
      automatic logic [1:0][31:0] _T_45 = {{Register_inst42}, {_T_1}};	// <stdin>:638:12, :649:12
      automatic logic [1:0][31:0] _T_46 = {{Register_inst43}, {_T_1}};	// <stdin>:653:12, :664:12
      automatic logic [1:0][31:0] _T_47 = {{Register_inst44}, {_T_1}};	// <stdin>:668:12, :679:12
      automatic logic [1:0][31:0] _T_48 = {{Register_inst45}, {_T_1}};	// <stdin>:683:12, :694:12
      automatic logic [1:0][31:0] _T_49 = {{Register_inst46}, {_T_1}};	// <stdin>:698:12, :709:12
      automatic logic [1:0][31:0] _T_50 = {{Register_inst47}, {_T_1}};	// <stdin>:713:12, :724:12
      automatic logic [1:0][31:0] _T_51 = {{Register_inst48}, {_T_1}};	// <stdin>:728:12, :739:12
      automatic logic [1:0][31:0] _T_52 = {{Register_inst49}, {_T_1}};	// <stdin>:743:12, :754:12
      automatic logic [1:0][31:0] _T_53 = {{Register_inst50}, {_T_1}};	// <stdin>:758:12, :769:12
      automatic logic [1:0][31:0] _T_54 = {{Register_inst51}, {_T_1}};	// <stdin>:773:12, :784:12
      automatic logic [1:0][31:0] _T_55 = {{Register_inst52}, {_T_1}};	// <stdin>:788:12, :799:12
      automatic logic [1:0][31:0] _T_56 = {{Register_inst53}, {_T_1}};	// <stdin>:803:12, :814:12
      automatic logic [1:0][31:0] _T_57 = {{Register_inst54}, {_T_1}};	// <stdin>:818:12, :829:12
      automatic logic [1:0][31:0] _T_58 = {{Register_inst55}, {_T_1}};	// <stdin>:833:12, :844:12
      automatic logic [1:0][31:0] _T_59 = {{Register_inst56}, {_T_1}};	// <stdin>:848:12, :859:12
      automatic logic [1:0][31:0] _T_60 = {{Register_inst57}, {_T_1}};	// <stdin>:863:12, :874:12
      automatic logic [1:0][31:0] _T_61 = {{Register_inst58}, {_T_1}};	// <stdin>:878:12, :889:12
      automatic logic [1:0][31:0] _T_62 = {{Register_inst59}, {_T_1}};	// <stdin>:893:12, :904:12
      automatic logic [1:0][31:0] _T_63 = {{Register_inst60}, {_T_1}};	// <stdin>:908:12, :919:12
      automatic logic [1:0][31:0] _T_64 = {{Register_inst61}, {_T_1}};	// <stdin>:923:12, :934:12
      automatic logic [1:0][31:0] _T_65 = {{Register_inst62}, {_T_1}};	// <stdin>:938:12, :949:12
      automatic logic [1:0][31:0] _T_66 = {{Register_inst63}, {_T_1}};	// <stdin>:953:12, :964:12
      automatic logic [1:0][31:0] _T_67 = {{Register_inst64}, {_T_1}};	// <stdin>:968:12, :979:12
      automatic logic [1:0][31:0] _T_68 = {{Register_inst65}, {_T_1}};	// <stdin>:983:12, :994:12
      automatic logic [1:0][31:0] _T_69 = {{Register_inst66}, {_T_1}};	// <stdin>:998:12, :1009:12
      automatic logic [1:0][31:0] _T_70 = {{Register_inst67}, {_T_1}};	// <stdin>:1013:12, :1024:12
      automatic logic [1:0][31:0] _T_71 = {{Register_inst68}, {_T_1}};	// <stdin>:1028:12, :1039:12
      automatic logic [1:0][31:0] _T_72 = {{Register_inst69}, {_T_1}};	// <stdin>:1043:12, :1054:12
      automatic logic [1:0][31:0] _T_73 = {{Register_inst70}, {_T_1}};	// <stdin>:1058:12, :1069:12
      automatic logic [1:0][31:0] _T_74 = {{Register_inst71}, {_T_1}};	// <stdin>:1073:12, :1084:12
      automatic logic [1:0][31:0] _T_75 = {{Register_inst72}, {_T_1}};	// <stdin>:1088:12, :1099:12
      automatic logic [1:0][31:0] _T_76 = {{Register_inst73}, {_T_1}};	// <stdin>:1103:12, :1114:12
      automatic logic [1:0][31:0] _T_77 = {{Register_inst74}, {_T_1}};	// <stdin>:1118:12, :1129:12
      automatic logic [1:0][31:0] _T_78 = {{Register_inst75}, {_T_1}};	// <stdin>:1133:12, :1144:12
      automatic logic [1:0][31:0] _T_79 = {{Register_inst76}, {_T_1}};	// <stdin>:1148:12, :1159:12
      automatic logic [1:0][31:0] _T_80 = {{Register_inst77}, {_T_1}};	// <stdin>:1163:12, :1174:12
      automatic logic [1:0][31:0] _T_81 = {{Register_inst78}, {_T_1}};	// <stdin>:1178:12, :1189:12
      automatic logic [1:0][31:0] _T_82 = {{Register_inst79}, {_T_1}};	// <stdin>:1193:12, :1204:12
      automatic logic [1:0][31:0] _T_83 = {{Register_inst80}, {_T_1}};	// <stdin>:1208:12, :1219:12
      automatic logic [1:0][31:0] _T_84 = {{Register_inst81}, {_T_1}};	// <stdin>:1223:12, :1234:12
      automatic logic [1:0][31:0] _T_85 = {{Register_inst82}, {_T_1}};	// <stdin>:1238:12, :1249:12
      automatic logic [1:0][31:0] _T_86 = {{Register_inst83}, {_T_1}};	// <stdin>:1253:12, :1264:12
      automatic logic [1:0][31:0] _T_87 = {{Register_inst84}, {_T_1}};	// <stdin>:1268:12, :1279:12
      automatic logic [1:0][31:0] _T_88 = {{Register_inst85}, {_T_1}};	// <stdin>:1283:12, :1294:12
      automatic logic [1:0][31:0] _T_89 = {{Register_inst86}, {_T_1}};	// <stdin>:1298:12, :1309:12
      automatic logic [1:0][31:0] _T_90 = {{Register_inst87}, {_T_1}};	// <stdin>:1313:12, :1324:12
      automatic logic [1:0][31:0] _T_91 = {{Register_inst88}, {_T_1}};	// <stdin>:1328:12, :1339:12
      automatic logic [1:0][31:0] _T_92 = {{Register_inst89}, {_T_1}};	// <stdin>:1343:12, :1354:12
      automatic logic [1:0][31:0] _T_93 = {{Register_inst90}, {_T_1}};	// <stdin>:1358:12, :1369:12
      automatic logic [1:0][31:0] _T_94 = {{Register_inst91}, {_T_1}};	// <stdin>:1373:12, :1384:12
      automatic logic [1:0][31:0] _T_95 = {{Register_inst92}, {_T_1}};	// <stdin>:1388:12, :1399:12
      automatic logic [1:0][31:0] _T_96 = {{Register_inst93}, {_T_1}};	// <stdin>:1403:12, :1414:12
      automatic logic [1:0][31:0] _T_97 = {{Register_inst94}, {_T_1}};	// <stdin>:1418:12, :1429:12
      automatic logic [1:0][31:0] _T_98 = {{Register_inst95}, {_T_1}};	// <stdin>:1433:12, :1444:12
      automatic logic [1:0][31:0] _T_99 = {{Register_inst96}, {_T_1}};	// <stdin>:1448:12, :1459:12
      automatic logic [1:0][31:0] _T_100 = {{Register_inst97}, {_T_1}};	// <stdin>:1463:12, :1474:12
      automatic logic [1:0][31:0] _T_101 = {{Register_inst98}, {_T_1}};	// <stdin>:1478:12, :1489:12
      automatic logic [1:0][31:0] _T_102 = {{Register_inst99}, {_T_1}};	// <stdin>:1493:12, :1504:12
      automatic logic [1:0][31:0] _T_103 = {{Register_inst100}, {_T_1}};	// <stdin>:1508:12, :1519:12
      automatic logic [1:0][31:0] _T_104 = {{Register_inst101}, {_T_1}};	// <stdin>:1523:12, :1534:12
      automatic logic [1:0][31:0] _T_105 = {{Register_inst102}, {_T_1}};	// <stdin>:1538:12, :1549:12
      automatic logic [1:0][31:0] _T_106 = {{Register_inst103}, {_T_1}};	// <stdin>:1553:12, :1564:12
      automatic logic [1:0][31:0] _T_107 = {{Register_inst104}, {_T_1}};	// <stdin>:1568:12, :1579:12
      automatic logic [1:0][31:0] _T_108 = {{Register_inst105}, {_T_1}};	// <stdin>:1583:12, :1594:12
      automatic logic [1:0][31:0] _T_109 = {{Register_inst106}, {_T_1}};	// <stdin>:1598:12, :1609:12
      automatic logic [1:0][31:0] _T_110 = {{Register_inst107}, {_T_1}};	// <stdin>:1613:12, :1624:12
      automatic logic [1:0][31:0] _T_111 = {{Register_inst108}, {_T_1}};	// <stdin>:1628:12, :1639:12
      automatic logic [1:0][31:0] _T_112 = {{Register_inst109}, {_T_1}};	// <stdin>:1643:12, :1654:12
      automatic logic [1:0][31:0] _T_113 = {{Register_inst110}, {_T_1}};	// <stdin>:1658:12, :1669:12
      automatic logic [1:0][31:0] _T_114 = {{Register_inst111}, {_T_1}};	// <stdin>:1673:12, :1684:12
      automatic logic [1:0][31:0] _T_115 = {{Register_inst112}, {_T_1}};	// <stdin>:1688:12, :1699:12
      automatic logic [1:0][31:0] _T_116 = {{Register_inst113}, {_T_1}};	// <stdin>:1703:12, :1714:12
      automatic logic [1:0][31:0] _T_117 = {{Register_inst114}, {_T_1}};	// <stdin>:1718:12, :1729:12
      automatic logic [1:0][31:0] _T_118 = {{Register_inst115}, {_T_1}};	// <stdin>:1733:12, :1744:12
      automatic logic [1:0][31:0] _T_119 = {{Register_inst116}, {_T_1}};	// <stdin>:1748:12, :1759:12
      automatic logic [1:0][31:0] _T_120 = {{Register_inst117}, {_T_1}};	// <stdin>:1763:12, :1774:12
      automatic logic [1:0][31:0] _T_121 = {{Register_inst118}, {_T_1}};	// <stdin>:1778:12, :1789:12
      automatic logic [1:0][31:0] _T_122 = {{Register_inst119}, {_T_1}};	// <stdin>:1793:12, :1804:12
      automatic logic [1:0][31:0] _T_123 = {{Register_inst120}, {_T_1}};	// <stdin>:1808:12, :1819:12
      automatic logic [1:0][31:0] _T_124 = {{Register_inst121}, {_T_1}};	// <stdin>:1823:12, :1834:12
      automatic logic [1:0][31:0] _T_125 = {{Register_inst122}, {_T_1}};	// <stdin>:1838:12, :1849:12
      automatic logic [1:0][31:0] _T_126 = {{Register_inst123}, {_T_1}};	// <stdin>:1853:12, :1864:12
      automatic logic [1:0][31:0] _T_127 = {{Register_inst124}, {_T_1}};	// <stdin>:1868:12, :1879:12
      automatic logic [1:0][31:0] _T_128 = {{Register_inst125}, {_T_1}};	// <stdin>:1883:12, :1894:12
      automatic logic [1:0][31:0] _T_129 = {{Register_inst126}, {_T_1}};	// <stdin>:1898:12, :1909:12
      automatic logic [1:0][31:0] _T_130 = {{Register_inst127}, {_T_1}};	// <stdin>:1913:12, :1924:12
      automatic logic [1:0][31:0] _T_131 = {{Register_inst128}, {_T_1}};	// <stdin>:1928:12, :1939:12
      automatic logic [1:0][31:0] _T_132 = {{Register_inst129}, {_T_1}};	// <stdin>:1943:12, :1954:12
      automatic logic [1:0][31:0] _T_133 = {{Register_inst130}, {_T_1}};	// <stdin>:1958:12, :1969:12
      automatic logic [1:0][31:0] _T_134 = {{Register_inst131}, {_T_1}};	// <stdin>:1973:12, :1984:12
      automatic logic [1:0][31:0] _T_135 = {{Register_inst132}, {_T_1}};	// <stdin>:1988:12, :1999:12
      automatic logic [1:0][31:0] _T_136 = {{Register_inst133}, {_T_1}};	// <stdin>:2003:12, :2014:12
      automatic logic [1:0][31:0] _T_137 = {{Register_inst134}, {_T_1}};	// <stdin>:2018:12, :2029:12
      automatic logic [1:0][31:0] _T_138 = {{Register_inst135}, {_T_1}};	// <stdin>:2033:12, :2044:12
      automatic logic [1:0][31:0] _T_139 = {{Register_inst136}, {_T_1}};	// <stdin>:2048:12, :2059:12
      automatic logic [1:0][31:0] _T_140 = {{Register_inst137}, {_T_1}};	// <stdin>:2063:12, :2074:12
      automatic logic [1:0][31:0] _T_141 = {{Register_inst138}, {_T_1}};	// <stdin>:2078:12, :2089:12
      automatic logic [1:0][31:0] _T_142 = {{Register_inst139}, {_T_1}};	// <stdin>:2093:12, :2104:12
      automatic logic [1:0][31:0] _T_143 = {{Register_inst140}, {_T_1}};	// <stdin>:2108:12, :2119:12
      automatic logic [1:0][31:0] _T_144 = {{Register_inst141}, {_T_1}};	// <stdin>:2123:12, :2134:12
      automatic logic [1:0][31:0] _T_145 = {{Register_inst142}, {_T_1}};	// <stdin>:2138:13, :2149:13
      automatic logic [1:0][31:0] _T_146 = {{Register_inst143}, {_T_1}};	// <stdin>:2153:13, :2164:13
      automatic logic [1:0][31:0] _T_147 = {{Register_inst144}, {_T_1}};	// <stdin>:2168:13, :2179:13
      automatic logic [1:0][31:0] _T_148 = {{Register_inst145}, {_T_1}};	// <stdin>:2183:13, :2194:13
      automatic logic [1:0][31:0] _T_149 = {{Register_inst146}, {_T_1}};	// <stdin>:2198:13, :2209:13
      automatic logic [1:0][31:0] _T_150 = {{Register_inst147}, {_T_1}};	// <stdin>:2213:13, :2224:13
      automatic logic [1:0][31:0] _T_151 = {{Register_inst148}, {_T_1}};	// <stdin>:2228:13, :2239:13
      automatic logic [1:0][31:0] _T_152 = {{Register_inst149}, {_T_1}};	// <stdin>:2243:13, :2254:13
      automatic logic [1:0][31:0] _T_153 = {{Register_inst150}, {_T_1}};	// <stdin>:2258:13, :2269:13
      automatic logic [1:0][31:0] _T_154 = {{Register_inst151}, {_T_1}};	// <stdin>:2273:13, :2284:13
      automatic logic [1:0][31:0] _T_155 = {{Register_inst152}, {_T_1}};	// <stdin>:2288:13, :2299:13
      automatic logic [1:0][31:0] _T_156 = {{Register_inst153}, {_T_1}};	// <stdin>:2303:13, :2314:13
      automatic logic [1:0][31:0] _T_157 = {{Register_inst154}, {_T_1}};	// <stdin>:2318:13, :2329:13
      automatic logic [1:0][31:0] _T_158 = {{Register_inst155}, {_T_1}};	// <stdin>:2333:13, :2344:13
      automatic logic [1:0][31:0] _T_159 = {{Register_inst156}, {_T_1}};	// <stdin>:2348:13, :2359:13
      automatic logic [1:0][31:0] _T_160 = {{Register_inst157}, {_T_1}};	// <stdin>:2363:13, :2374:13
      automatic logic [1:0][31:0] _T_161 = {{Register_inst158}, {_T_1}};	// <stdin>:2378:13, :2389:13
      automatic logic [1:0][31:0] _T_162 = {{Register_inst159}, {_T_1}};	// <stdin>:2393:13, :2404:13
      automatic logic [1:0][31:0] _T_163 = {{Register_inst160}, {_T_1}};	// <stdin>:2408:13, :2419:13
      automatic logic [1:0][31:0] _T_164 = {{Register_inst161}, {_T_1}};	// <stdin>:2423:13, :2434:13
      automatic logic [1:0][31:0] _T_165 = {{Register_inst162}, {_T_1}};	// <stdin>:2438:13, :2449:13
      automatic logic [1:0][31:0] _T_166 = {{Register_inst163}, {_T_1}};	// <stdin>:2453:13, :2464:13
      automatic logic [1:0][31:0] _T_167 = {{Register_inst164}, {_T_1}};	// <stdin>:2468:13, :2479:13
      automatic logic [1:0][31:0] _T_168 = {{Register_inst165}, {_T_1}};	// <stdin>:2483:13, :2494:13
      automatic logic [1:0][31:0] _T_169 = {{Register_inst166}, {_T_1}};	// <stdin>:2498:13, :2509:13
      automatic logic [1:0][31:0] _T_170 = {{Register_inst167}, {_T_1}};	// <stdin>:2513:13, :2524:13
      automatic logic [1:0][31:0] _T_171 = {{Register_inst168}, {_T_1}};	// <stdin>:2528:13, :2539:13
      automatic logic [1:0][31:0] _T_172 = {{Register_inst169}, {_T_1}};	// <stdin>:2543:13, :2554:13
      automatic logic [1:0][31:0] _T_173 = {{Register_inst170}, {_T_1}};	// <stdin>:2558:13, :2569:13
      automatic logic [1:0][31:0] _T_174 = {{Register_inst171}, {_T_1}};	// <stdin>:2573:13, :2584:13
      automatic logic [1:0][31:0] _T_175 = {{Register_inst172}, {_T_1}};	// <stdin>:2588:13, :2599:13
      automatic logic [1:0][31:0] _T_176 = {{Register_inst173}, {_T_1}};	// <stdin>:2603:13, :2614:13
      automatic logic [1:0][31:0] _T_177 = {{Register_inst174}, {_T_1}};	// <stdin>:2618:13, :2629:13
      automatic logic [1:0][31:0] _T_178 = {{Register_inst175}, {_T_1}};	// <stdin>:2633:13, :2644:13
      automatic logic [1:0][31:0] _T_179 = {{Register_inst176}, {_T_1}};	// <stdin>:2648:13, :2659:13
      automatic logic [1:0][31:0] _T_180 = {{Register_inst177}, {_T_1}};	// <stdin>:2663:13, :2674:13
      automatic logic [1:0][31:0] _T_181 = {{Register_inst178}, {_T_1}};	// <stdin>:2678:13, :2689:13
      automatic logic [1:0][31:0] _T_182 = {{Register_inst179}, {_T_1}};	// <stdin>:2693:13, :2704:13
      automatic logic [1:0][31:0] _T_183 = {{Register_inst180}, {_T_1}};	// <stdin>:2708:13, :2719:13
      automatic logic [1:0][31:0] _T_184 = {{Register_inst181}, {_T_1}};	// <stdin>:2723:13, :2734:13
      automatic logic [1:0][31:0] _T_185 = {{Register_inst182}, {_T_1}};	// <stdin>:2738:13, :2749:13
      automatic logic [1:0][31:0] _T_186 = {{Register_inst183}, {_T_1}};	// <stdin>:2753:13, :2764:13
      automatic logic [1:0][31:0] _T_187 = {{Register_inst184}, {_T_1}};	// <stdin>:2768:13, :2779:13
      automatic logic [1:0][31:0] _T_188 = {{Register_inst185}, {_T_1}};	// <stdin>:2783:13, :2794:13
      automatic logic [1:0][31:0] _T_189 = {{Register_inst186}, {_T_1}};	// <stdin>:2798:13, :2809:13
      automatic logic [1:0][31:0] _T_190 = {{Register_inst187}, {_T_1}};	// <stdin>:2813:13, :2824:13
      automatic logic [1:0][31:0] _T_191 = {{Register_inst188}, {_T_1}};	// <stdin>:2828:13, :2839:13
      automatic logic [1:0][31:0] _T_192 = {{Register_inst189}, {_T_1}};	// <stdin>:2843:13, :2854:13
      automatic logic [1:0][31:0] _T_193 = {{Register_inst190}, {_T_1}};	// <stdin>:2858:13, :2869:13
      automatic logic [1:0][31:0] _T_194 = {{Register_inst191}, {_T_1}};	// <stdin>:2873:13, :2884:13
      automatic logic [1:0][31:0] _T_195 = {{Register_inst192}, {_T_1}};	// <stdin>:2888:13, :2899:13
      automatic logic [1:0][31:0] _T_196 = {{Register_inst193}, {_T_1}};	// <stdin>:2903:13, :2914:13
      automatic logic [1:0][31:0] _T_197 = {{Register_inst194}, {_T_1}};	// <stdin>:2918:13, :2929:13
      automatic logic [1:0][31:0] _T_198 = {{Register_inst195}, {_T_1}};	// <stdin>:2933:13, :2944:13
      automatic logic [1:0][31:0] _T_199 = {{Register_inst196}, {_T_1}};	// <stdin>:2948:13, :2959:13
      automatic logic [1:0][31:0] _T_200 = {{Register_inst197}, {_T_1}};	// <stdin>:2963:13, :2974:13
      automatic logic [1:0][31:0] _T_201 = {{Register_inst198}, {_T_1}};	// <stdin>:2978:13, :2989:13
      automatic logic [1:0][31:0] _T_202 = {{Register_inst199}, {_T_1}};	// <stdin>:2993:13, :3004:13
      automatic logic [1:0][31:0] _T_203 = {{Register_inst200}, {_T_1}};	// <stdin>:3008:13, :3019:13
      automatic logic [1:0][31:0] _T_204 = {{Register_inst201}, {_T_1}};	// <stdin>:3023:13, :3034:13
      automatic logic [1:0][31:0] _T_205 = {{Register_inst202}, {_T_1}};	// <stdin>:3038:13, :3049:13
      automatic logic [1:0][31:0] _T_206 = {{Register_inst203}, {_T_1}};	// <stdin>:3053:13, :3064:13
      automatic logic [1:0][31:0] _T_207 = {{Register_inst204}, {_T_1}};	// <stdin>:3068:13, :3079:13
      automatic logic [1:0][31:0] _T_208 = {{Register_inst205}, {_T_1}};	// <stdin>:3083:13, :3094:13
      automatic logic [1:0][31:0] _T_209 = {{Register_inst206}, {_T_1}};	// <stdin>:3098:13, :3109:13
      automatic logic [1:0][31:0] _T_210 = {{Register_inst207}, {_T_1}};	// <stdin>:3113:13, :3124:13
      automatic logic [1:0][31:0] _T_211 = {{Register_inst208}, {_T_1}};	// <stdin>:3128:13, :3139:13
      automatic logic [1:0][31:0] _T_212 = {{Register_inst209}, {_T_1}};	// <stdin>:3143:13, :3154:13
      automatic logic [1:0][31:0] _T_213 = {{Register_inst210}, {_T_1}};	// <stdin>:3158:13, :3169:13
      automatic logic [1:0][31:0] _T_214 = {{Register_inst211}, {_T_1}};	// <stdin>:3173:13, :3184:13
      automatic logic [1:0][31:0] _T_215 = {{Register_inst212}, {_T_1}};	// <stdin>:3188:13, :3199:13
      automatic logic [1:0][31:0] _T_216 = {{Register_inst213}, {_T_1}};	// <stdin>:3203:13, :3214:13
      automatic logic [1:0][31:0] _T_217 = {{Register_inst214}, {_T_1}};	// <stdin>:3218:13, :3229:13
      automatic logic [1:0][31:0] _T_218 = {{Register_inst215}, {_T_1}};	// <stdin>:3233:13, :3244:13
      automatic logic [1:0][31:0] _T_219 = {{Register_inst216}, {_T_1}};	// <stdin>:3248:13, :3259:13
      automatic logic [1:0][31:0] _T_220 = {{Register_inst217}, {_T_1}};	// <stdin>:3263:13, :3274:13
      automatic logic [1:0][31:0] _T_221 = {{Register_inst218}, {_T_1}};	// <stdin>:3278:13, :3289:13
      automatic logic [1:0][31:0] _T_222 = {{Register_inst219}, {_T_1}};	// <stdin>:3293:13, :3304:13
      automatic logic [1:0][31:0] _T_223 = {{Register_inst220}, {_T_1}};	// <stdin>:3308:13, :3319:13
      automatic logic [1:0][31:0] _T_224 = {{Register_inst221}, {_T_1}};	// <stdin>:3323:13, :3334:13
      automatic logic [1:0][31:0] _T_225 = {{Register_inst222}, {_T_1}};	// <stdin>:3338:13, :3349:13
      automatic logic [1:0][31:0] _T_226 = {{Register_inst223}, {_T_1}};	// <stdin>:3353:13, :3364:13
      automatic logic [1:0][31:0] _T_227 = {{Register_inst224}, {_T_1}};	// <stdin>:3368:13, :3379:13
      automatic logic [1:0][31:0] _T_228 = {{Register_inst225}, {_T_1}};	// <stdin>:3383:13, :3394:13
      automatic logic [1:0][31:0] _T_229 = {{Register_inst226}, {_T_1}};	// <stdin>:3398:13, :3409:13
      automatic logic [1:0][31:0] _T_230 = {{Register_inst227}, {_T_1}};	// <stdin>:3413:13, :3424:13
      automatic logic [1:0][31:0] _T_231 = {{Register_inst228}, {_T_1}};	// <stdin>:3428:13, :3439:13
      automatic logic [1:0][31:0] _T_232 = {{Register_inst229}, {_T_1}};	// <stdin>:3443:13, :3454:13
      automatic logic [1:0][31:0] _T_233 = {{Register_inst230}, {_T_1}};	// <stdin>:3458:13, :3469:13
      automatic logic [1:0][31:0] _T_234 = {{Register_inst231}, {_T_1}};	// <stdin>:3473:13, :3484:13
      automatic logic [1:0][31:0] _T_235 = {{Register_inst232}, {_T_1}};	// <stdin>:3488:13, :3499:13
      automatic logic [1:0][31:0] _T_236 = {{Register_inst233}, {_T_1}};	// <stdin>:3503:13, :3514:13
      automatic logic [1:0][31:0] _T_237 = {{Register_inst234}, {_T_1}};	// <stdin>:3518:13, :3529:13
      automatic logic [1:0][31:0] _T_238 = {{Register_inst235}, {_T_1}};	// <stdin>:3533:13, :3544:13
      automatic logic [1:0][31:0] _T_239 = {{Register_inst236}, {_T_1}};	// <stdin>:3548:13, :3559:13
      automatic logic [1:0][31:0] _T_240 = {{Register_inst237}, {_T_1}};	// <stdin>:3563:13, :3574:13
      automatic logic [1:0][31:0] _T_241 = {{Register_inst238}, {_T_1}};	// <stdin>:3578:13, :3589:13
      automatic logic [1:0][31:0] _T_242 = {{Register_inst239}, {_T_1}};	// <stdin>:3593:13, :3604:13
      automatic logic [1:0][31:0] _T_243 = {{Register_inst240}, {_T_1}};	// <stdin>:3608:13, :3619:13
      automatic logic [1:0][31:0] _T_244 = {{Register_inst241}, {_T_1}};	// <stdin>:3623:13, :3634:13
      automatic logic [1:0][31:0] _T_245 = {{Register_inst242}, {_T_1}};	// <stdin>:3638:13, :3649:13
      automatic logic [1:0][31:0] _T_246 = {{Register_inst243}, {_T_1}};	// <stdin>:3653:13, :3664:13
      automatic logic [1:0][31:0] _T_247 = {{Register_inst244}, {_T_1}};	// <stdin>:3668:13, :3679:13
      automatic logic [1:0][31:0] _T_248 = {{Register_inst245}, {_T_1}};	// <stdin>:3683:13, :3694:13
      automatic logic [1:0][31:0] _T_249 = {{Register_inst246}, {_T_1}};	// <stdin>:3698:13, :3709:13
      automatic logic [1:0][31:0] _T_250 = {{Register_inst247}, {_T_1}};	// <stdin>:3713:13, :3724:13
      automatic logic [1:0][31:0] _T_251 = {{Register_inst248}, {_T_1}};	// <stdin>:3728:13, :3739:13
      automatic logic [1:0][31:0] _T_252 = {{Register_inst249}, {_T_1}};	// <stdin>:3743:13, :3754:13
      automatic logic [1:0][31:0] _T_253 = {{Register_inst250}, {_T_1}};	// <stdin>:3758:13, :3769:13
      automatic logic [1:0][31:0] _T_254 = {{Register_inst251}, {_T_1}};	// <stdin>:3773:13, :3784:13
      automatic logic [1:0][31:0] _T_255 = {{Register_inst252}, {_T_1}};	// <stdin>:3788:13, :3799:13
      automatic logic [1:0][31:0] _T_256 = {{Register_inst253}, {_T_1}};	// <stdin>:3803:13, :3814:13
      automatic logic [1:0][31:0] _T_257 = {{Register_inst254}, {_T_1}};	// <stdin>:3818:13, :3829:13
      automatic logic [1:0][31:0] _T_258 = {{Register_inst255}, {_T_1}};	// <stdin>:3833:13, :3844:13

      Register_inst0 <= _T_3[_T_2 == 8'h0 & write_0_en];	// <stdin>:4:10, :5:10, :6:10, :8:10, :11:9
      Register_inst1 <= _T_4[_T_2 == 8'h1 & write_0_en];	// <stdin>:20:11, :21:11, :22:11, :24:11, :27:9
      Register_inst2 <= _T_5[_T_2 == 8'h2 & write_0_en];	// <stdin>:35:11, :36:11, :37:11, :39:11, :42:9
      Register_inst3 <= _T_6[_T_2 == 8'h3 & write_0_en];	// <stdin>:50:11, :51:11, :52:11, :54:11, :57:9
      Register_inst4 <= _T_7[_T_2 == 8'h4 & write_0_en];	// <stdin>:65:11, :66:11, :67:11, :69:11, :72:9
      Register_inst5 <= _T_8[_T_2 == 8'h5 & write_0_en];	// <stdin>:80:11, :81:11, :82:11, :84:11, :87:9
      Register_inst6 <= _T_9[_T_2 == 8'h6 & write_0_en];	// <stdin>:95:11, :96:11, :97:11, :99:11, :102:9
      Register_inst7 <= _T_10[_T_2 == 8'h7 & write_0_en];	// <stdin>:110:11, :111:11, :112:11, :114:11, :117:9
      Register_inst8 <= _T_11[_T_2 == 8'h8 & write_0_en];	// <stdin>:125:11, :126:11, :127:11, :129:11, :132:9
      Register_inst9 <= _T_12[_T_2 == 8'h9 & write_0_en];	// <stdin>:140:11, :141:11, :142:11, :144:11, :147:9
      Register_inst10 <= _T_13[_T_2 == 8'hA & write_0_en];	// <stdin>:155:11, :156:11, :157:11, :159:11, :162:9
      Register_inst11 <= _T_14[_T_2 == 8'hB & write_0_en];	// <stdin>:170:11, :171:11, :172:11, :174:11, :177:9
      Register_inst12 <= _T_15[_T_2 == 8'hC & write_0_en];	// <stdin>:185:11, :186:11, :187:11, :189:11, :192:9
      Register_inst13 <= _T_16[_T_2 == 8'hD & write_0_en];	// <stdin>:200:11, :201:11, :202:11, :204:11, :207:9
      Register_inst14 <= _T_17[_T_2 == 8'hE & write_0_en];	// <stdin>:215:12, :216:12, :217:12, :219:12, :222:9
      Register_inst15 <= _T_18[_T_2 == 8'hF & write_0_en];	// <stdin>:230:12, :231:12, :232:12, :234:12, :237:9
      Register_inst16 <= _T_19[_T_2 == 8'h10 & write_0_en];	// <stdin>:245:12, :246:12, :247:12, :249:12, :252:9
      Register_inst17 <= _T_20[_T_2 == 8'h11 & write_0_en];	// <stdin>:260:12, :261:12, :262:12, :264:12, :267:9
      Register_inst18 <= _T_21[_T_2 == 8'h12 & write_0_en];	// <stdin>:275:12, :276:12, :277:12, :279:12, :282:9
      Register_inst19 <= _T_22[_T_2 == 8'h13 & write_0_en];	// <stdin>:290:12, :291:12, :292:12, :294:12, :297:9
      Register_inst20 <= _T_23[_T_2 == 8'h14 & write_0_en];	// <stdin>:305:12, :306:12, :307:12, :309:12, :312:9
      Register_inst21 <= _T_24[_T_2 == 8'h15 & write_0_en];	// <stdin>:320:12, :321:12, :322:12, :324:12, :327:9
      Register_inst22 <= _T_25[_T_2 == 8'h16 & write_0_en];	// <stdin>:335:12, :336:12, :337:12, :339:12, :342:9
      Register_inst23 <= _T_26[_T_2 == 8'h17 & write_0_en];	// <stdin>:350:12, :351:12, :352:12, :354:12, :357:9
      Register_inst24 <= _T_27[_T_2 == 8'h18 & write_0_en];	// <stdin>:365:12, :366:12, :367:12, :369:12, :372:9
      Register_inst25 <= _T_28[_T_2 == 8'h19 & write_0_en];	// <stdin>:380:12, :381:12, :382:12, :384:12, :387:9
      Register_inst26 <= _T_29[_T_2 == 8'h1A & write_0_en];	// <stdin>:395:12, :396:12, :397:12, :399:12, :402:9
      Register_inst27 <= _T_30[_T_2 == 8'h1B & write_0_en];	// <stdin>:410:12, :411:12, :412:12, :414:12, :417:9
      Register_inst28 <= _T_31[_T_2 == 8'h1C & write_0_en];	// <stdin>:425:12, :426:12, :427:12, :429:12, :432:9
      Register_inst29 <= _T_32[_T_2 == 8'h1D & write_0_en];	// <stdin>:440:12, :441:12, :442:12, :444:12, :447:9
      Register_inst30 <= _T_33[_T_2 == 8'h1E & write_0_en];	// <stdin>:455:12, :456:12, :457:12, :459:12, :462:9
      Register_inst31 <= _T_34[_T_2 == 8'h1F & write_0_en];	// <stdin>:470:12, :471:12, :472:12, :474:12, :477:9
      Register_inst32 <= _T_35[_T_2 == 8'h20 & write_0_en];	// <stdin>:485:12, :486:12, :487:12, :489:12, :492:9
      Register_inst33 <= _T_36[_T_2 == 8'h21 & write_0_en];	// <stdin>:500:12, :501:12, :502:12, :504:12, :507:9
      Register_inst34 <= _T_37[_T_2 == 8'h22 & write_0_en];	// <stdin>:515:12, :516:12, :517:12, :519:12, :522:9
      Register_inst35 <= _T_38[_T_2 == 8'h23 & write_0_en];	// <stdin>:530:12, :531:12, :532:12, :534:12, :537:9
      Register_inst36 <= _T_39[_T_2 == 8'h24 & write_0_en];	// <stdin>:545:12, :546:12, :547:12, :549:12, :552:9
      Register_inst37 <= _T_40[_T_2 == 8'h25 & write_0_en];	// <stdin>:560:12, :561:12, :562:12, :564:12, :567:9
      Register_inst38 <= _T_41[_T_2 == 8'h26 & write_0_en];	// <stdin>:575:12, :576:12, :577:12, :579:12, :582:9
      Register_inst39 <= _T_42[_T_2 == 8'h27 & write_0_en];	// <stdin>:590:12, :591:12, :592:12, :594:12, :597:9
      Register_inst40 <= _T_43[_T_2 == 8'h28 & write_0_en];	// <stdin>:605:12, :606:12, :607:12, :609:12, :612:9
      Register_inst41 <= _T_44[_T_2 == 8'h29 & write_0_en];	// <stdin>:620:12, :621:12, :622:12, :624:12, :627:9
      Register_inst42 <= _T_45[_T_2 == 8'h2A & write_0_en];	// <stdin>:635:12, :636:12, :637:12, :639:12, :642:9
      Register_inst43 <= _T_46[_T_2 == 8'h2B & write_0_en];	// <stdin>:650:12, :651:12, :652:12, :654:12, :657:9
      Register_inst44 <= _T_47[_T_2 == 8'h2C & write_0_en];	// <stdin>:665:12, :666:12, :667:12, :669:12, :672:9
      Register_inst45 <= _T_48[_T_2 == 8'h2D & write_0_en];	// <stdin>:680:12, :681:12, :682:12, :684:12, :687:9
      Register_inst46 <= _T_49[_T_2 == 8'h2E & write_0_en];	// <stdin>:695:12, :696:12, :697:12, :699:12, :702:9
      Register_inst47 <= _T_50[_T_2 == 8'h2F & write_0_en];	// <stdin>:710:12, :711:12, :712:12, :714:12, :717:9
      Register_inst48 <= _T_51[_T_2 == 8'h30 & write_0_en];	// <stdin>:725:12, :726:12, :727:12, :729:12, :732:9
      Register_inst49 <= _T_52[_T_2 == 8'h31 & write_0_en];	// <stdin>:740:12, :741:12, :742:12, :744:12, :747:9
      Register_inst50 <= _T_53[_T_2 == 8'h32 & write_0_en];	// <stdin>:755:12, :756:12, :757:12, :759:12, :762:9
      Register_inst51 <= _T_54[_T_2 == 8'h33 & write_0_en];	// <stdin>:770:12, :771:12, :772:12, :774:12, :777:9
      Register_inst52 <= _T_55[_T_2 == 8'h34 & write_0_en];	// <stdin>:785:12, :786:12, :787:12, :789:12, :792:9
      Register_inst53 <= _T_56[_T_2 == 8'h35 & write_0_en];	// <stdin>:800:12, :801:12, :802:12, :804:12, :807:9
      Register_inst54 <= _T_57[_T_2 == 8'h36 & write_0_en];	// <stdin>:815:12, :816:12, :817:12, :819:12, :822:9
      Register_inst55 <= _T_58[_T_2 == 8'h37 & write_0_en];	// <stdin>:830:12, :831:12, :832:12, :834:12, :837:9
      Register_inst56 <= _T_59[_T_2 == 8'h38 & write_0_en];	// <stdin>:845:12, :846:12, :847:12, :849:12, :852:9
      Register_inst57 <= _T_60[_T_2 == 8'h39 & write_0_en];	// <stdin>:860:12, :861:12, :862:12, :864:12, :867:9
      Register_inst58 <= _T_61[_T_2 == 8'h3A & write_0_en];	// <stdin>:875:12, :876:12, :877:12, :879:12, :882:9
      Register_inst59 <= _T_62[_T_2 == 8'h3B & write_0_en];	// <stdin>:890:12, :891:12, :892:12, :894:12, :897:9
      Register_inst60 <= _T_63[_T_2 == 8'h3C & write_0_en];	// <stdin>:905:12, :906:12, :907:12, :909:12, :912:9
      Register_inst61 <= _T_64[_T_2 == 8'h3D & write_0_en];	// <stdin>:920:12, :921:12, :922:12, :924:12, :927:9
      Register_inst62 <= _T_65[_T_2 == 8'h3E & write_0_en];	// <stdin>:935:12, :936:12, :937:12, :939:12, :942:9
      Register_inst63 <= _T_66[_T_2 == 8'h3F & write_0_en];	// <stdin>:950:12, :951:12, :952:12, :954:12, :957:9
      Register_inst64 <= _T_67[_T_2 == 8'h40 & write_0_en];	// <stdin>:965:12, :966:12, :967:12, :969:12, :972:9
      Register_inst65 <= _T_68[_T_2 == 8'h41 & write_0_en];	// <stdin>:980:12, :981:12, :982:12, :984:12, :987:9
      Register_inst66 <= _T_69[_T_2 == 8'h42 & write_0_en];	// <stdin>:995:12, :996:12, :997:12, :999:12, :1002:9
      Register_inst67 <= _T_70[_T_2 == 8'h43 & write_0_en];	// <stdin>:1010:12, :1011:12, :1012:12, :1014:12, :1017:9
      Register_inst68 <= _T_71[_T_2 == 8'h44 & write_0_en];	// <stdin>:1025:12, :1026:12, :1027:12, :1029:12, :1032:9
      Register_inst69 <= _T_72[_T_2 == 8'h45 & write_0_en];	// <stdin>:1040:12, :1041:12, :1042:12, :1044:12, :1047:9
      Register_inst70 <= _T_73[_T_2 == 8'h46 & write_0_en];	// <stdin>:1055:12, :1056:12, :1057:12, :1059:12, :1062:9
      Register_inst71 <= _T_74[_T_2 == 8'h47 & write_0_en];	// <stdin>:1070:12, :1071:12, :1072:12, :1074:12, :1077:9
      Register_inst72 <= _T_75[_T_2 == 8'h48 & write_0_en];	// <stdin>:1085:12, :1086:12, :1087:12, :1089:12, :1092:9
      Register_inst73 <= _T_76[_T_2 == 8'h49 & write_0_en];	// <stdin>:1100:12, :1101:12, :1102:12, :1104:12, :1107:9
      Register_inst74 <= _T_77[_T_2 == 8'h4A & write_0_en];	// <stdin>:1115:12, :1116:12, :1117:12, :1119:12, :1122:9
      Register_inst75 <= _T_78[_T_2 == 8'h4B & write_0_en];	// <stdin>:1130:12, :1131:12, :1132:12, :1134:12, :1137:9
      Register_inst76 <= _T_79[_T_2 == 8'h4C & write_0_en];	// <stdin>:1145:12, :1146:12, :1147:12, :1149:12, :1152:9
      Register_inst77 <= _T_80[_T_2 == 8'h4D & write_0_en];	// <stdin>:1160:12, :1161:12, :1162:12, :1164:12, :1167:9
      Register_inst78 <= _T_81[_T_2 == 8'h4E & write_0_en];	// <stdin>:1175:12, :1176:12, :1177:12, :1179:12, :1182:9
      Register_inst79 <= _T_82[_T_2 == 8'h4F & write_0_en];	// <stdin>:1190:12, :1191:12, :1192:12, :1194:12, :1197:9
      Register_inst80 <= _T_83[_T_2 == 8'h50 & write_0_en];	// <stdin>:1205:12, :1206:12, :1207:12, :1209:12, :1212:9
      Register_inst81 <= _T_84[_T_2 == 8'h51 & write_0_en];	// <stdin>:1220:12, :1221:12, :1222:12, :1224:12, :1227:9
      Register_inst82 <= _T_85[_T_2 == 8'h52 & write_0_en];	// <stdin>:1235:12, :1236:12, :1237:12, :1239:12, :1242:9
      Register_inst83 <= _T_86[_T_2 == 8'h53 & write_0_en];	// <stdin>:1250:12, :1251:12, :1252:12, :1254:12, :1257:9
      Register_inst84 <= _T_87[_T_2 == 8'h54 & write_0_en];	// <stdin>:1265:12, :1266:12, :1267:12, :1269:12, :1272:9
      Register_inst85 <= _T_88[_T_2 == 8'h55 & write_0_en];	// <stdin>:1280:12, :1281:12, :1282:12, :1284:12, :1287:9
      Register_inst86 <= _T_89[_T_2 == 8'h56 & write_0_en];	// <stdin>:1295:12, :1296:12, :1297:12, :1299:12, :1302:9
      Register_inst87 <= _T_90[_T_2 == 8'h57 & write_0_en];	// <stdin>:1310:12, :1311:12, :1312:12, :1314:12, :1317:9
      Register_inst88 <= _T_91[_T_2 == 8'h58 & write_0_en];	// <stdin>:1325:12, :1326:12, :1327:12, :1329:12, :1332:9
      Register_inst89 <= _T_92[_T_2 == 8'h59 & write_0_en];	// <stdin>:1340:12, :1341:12, :1342:12, :1344:12, :1347:9
      Register_inst90 <= _T_93[_T_2 == 8'h5A & write_0_en];	// <stdin>:1355:12, :1356:12, :1357:12, :1359:12, :1362:9
      Register_inst91 <= _T_94[_T_2 == 8'h5B & write_0_en];	// <stdin>:1370:12, :1371:12, :1372:12, :1374:12, :1377:9
      Register_inst92 <= _T_95[_T_2 == 8'h5C & write_0_en];	// <stdin>:1385:12, :1386:12, :1387:12, :1389:12, :1392:9
      Register_inst93 <= _T_96[_T_2 == 8'h5D & write_0_en];	// <stdin>:1400:12, :1401:12, :1402:12, :1404:12, :1407:9
      Register_inst94 <= _T_97[_T_2 == 8'h5E & write_0_en];	// <stdin>:1415:12, :1416:12, :1417:12, :1419:12, :1422:9
      Register_inst95 <= _T_98[_T_2 == 8'h5F & write_0_en];	// <stdin>:1430:12, :1431:12, :1432:12, :1434:12, :1437:9
      Register_inst96 <= _T_99[_T_2 == 8'h60 & write_0_en];	// <stdin>:1445:12, :1446:12, :1447:12, :1449:12, :1452:9
      Register_inst97 <= _T_100[_T_2 == 8'h61 & write_0_en];	// <stdin>:1460:12, :1461:12, :1462:12, :1464:12, :1467:9
      Register_inst98 <= _T_101[_T_2 == 8'h62 & write_0_en];	// <stdin>:1475:12, :1476:12, :1477:12, :1479:12, :1482:9
      Register_inst99 <= _T_102[_T_2 == 8'h63 & write_0_en];	// <stdin>:1490:12, :1491:12, :1492:12, :1494:12, :1497:9
      Register_inst100 <= _T_103[_T_2 == 8'h64 & write_0_en];	// <stdin>:1505:12, :1506:12, :1507:12, :1509:12, :1512:9
      Register_inst101 <= _T_104[_T_2 == 8'h65 & write_0_en];	// <stdin>:1520:12, :1521:12, :1522:12, :1524:12, :1527:9
      Register_inst102 <= _T_105[_T_2 == 8'h66 & write_0_en];	// <stdin>:1535:12, :1536:12, :1537:12, :1539:12, :1542:9
      Register_inst103 <= _T_106[_T_2 == 8'h67 & write_0_en];	// <stdin>:1550:12, :1551:12, :1552:12, :1554:12, :1557:9
      Register_inst104 <= _T_107[_T_2 == 8'h68 & write_0_en];	// <stdin>:1565:12, :1566:12, :1567:12, :1569:12, :1572:9
      Register_inst105 <= _T_108[_T_2 == 8'h69 & write_0_en];	// <stdin>:1580:12, :1581:12, :1582:12, :1584:12, :1587:9
      Register_inst106 <= _T_109[_T_2 == 8'h6A & write_0_en];	// <stdin>:1595:12, :1596:12, :1597:12, :1599:12, :1602:9
      Register_inst107 <= _T_110[_T_2 == 8'h6B & write_0_en];	// <stdin>:1610:12, :1611:12, :1612:12, :1614:12, :1617:9
      Register_inst108 <= _T_111[_T_2 == 8'h6C & write_0_en];	// <stdin>:1625:12, :1626:12, :1627:12, :1629:12, :1632:9
      Register_inst109 <= _T_112[_T_2 == 8'h6D & write_0_en];	// <stdin>:1640:12, :1641:12, :1642:12, :1644:12, :1647:9
      Register_inst110 <= _T_113[_T_2 == 8'h6E & write_0_en];	// <stdin>:1655:12, :1656:12, :1657:12, :1659:12, :1662:9
      Register_inst111 <= _T_114[_T_2 == 8'h6F & write_0_en];	// <stdin>:1670:12, :1671:12, :1672:12, :1674:12, :1677:9
      Register_inst112 <= _T_115[_T_2 == 8'h70 & write_0_en];	// <stdin>:1685:12, :1686:12, :1687:12, :1689:12, :1692:9
      Register_inst113 <= _T_116[_T_2 == 8'h71 & write_0_en];	// <stdin>:1700:12, :1701:12, :1702:12, :1704:12, :1707:9
      Register_inst114 <= _T_117[_T_2 == 8'h72 & write_0_en];	// <stdin>:1715:12, :1716:12, :1717:12, :1719:12, :1722:9
      Register_inst115 <= _T_118[_T_2 == 8'h73 & write_0_en];	// <stdin>:1730:12, :1731:12, :1732:12, :1734:12, :1737:9
      Register_inst116 <= _T_119[_T_2 == 8'h74 & write_0_en];	// <stdin>:1745:12, :1746:12, :1747:12, :1749:12, :1752:9
      Register_inst117 <= _T_120[_T_2 == 8'h75 & write_0_en];	// <stdin>:1760:12, :1761:12, :1762:12, :1764:12, :1767:9
      Register_inst118 <= _T_121[_T_2 == 8'h76 & write_0_en];	// <stdin>:1775:12, :1776:12, :1777:12, :1779:12, :1782:9
      Register_inst119 <= _T_122[_T_2 == 8'h77 & write_0_en];	// <stdin>:1790:12, :1791:12, :1792:12, :1794:12, :1797:9
      Register_inst120 <= _T_123[_T_2 == 8'h78 & write_0_en];	// <stdin>:1805:12, :1806:12, :1807:12, :1809:12, :1812:9
      Register_inst121 <= _T_124[_T_2 == 8'h79 & write_0_en];	// <stdin>:1820:12, :1821:12, :1822:12, :1824:12, :1827:9
      Register_inst122 <= _T_125[_T_2 == 8'h7A & write_0_en];	// <stdin>:1835:12, :1836:12, :1837:12, :1839:12, :1842:9
      Register_inst123 <= _T_126[_T_2 == 8'h7B & write_0_en];	// <stdin>:1850:12, :1851:12, :1852:12, :1854:12, :1857:9
      Register_inst124 <= _T_127[_T_2 == 8'h7C & write_0_en];	// <stdin>:1865:12, :1866:12, :1867:12, :1869:12, :1872:9
      Register_inst125 <= _T_128[_T_2 == 8'h7D & write_0_en];	// <stdin>:1880:12, :1881:12, :1882:12, :1884:12, :1887:9
      Register_inst126 <= _T_129[_T_2 == 8'h7E & write_0_en];	// <stdin>:1895:12, :1896:12, :1897:12, :1899:12, :1902:9
      Register_inst127 <= _T_130[_T_2 == 8'h7F & write_0_en];	// <stdin>:1910:12, :1911:12, :1912:12, :1914:12, :1917:9
      Register_inst128 <= _T_131[_T_2 == 8'h80 & write_0_en];	// <stdin>:1925:12, :1926:12, :1927:12, :1929:12, :1932:9
      Register_inst129 <= _T_132[_T_2 == 8'h81 & write_0_en];	// <stdin>:1940:12, :1941:12, :1942:12, :1944:12, :1947:9
      Register_inst130 <= _T_133[_T_2 == 8'h82 & write_0_en];	// <stdin>:1955:12, :1956:12, :1957:12, :1959:12, :1962:9
      Register_inst131 <= _T_134[_T_2 == 8'h83 & write_0_en];	// <stdin>:1970:12, :1971:12, :1972:12, :1974:12, :1977:9
      Register_inst132 <= _T_135[_T_2 == 8'h84 & write_0_en];	// <stdin>:1985:12, :1986:12, :1987:12, :1989:12, :1992:9
      Register_inst133 <= _T_136[_T_2 == 8'h85 & write_0_en];	// <stdin>:2000:12, :2001:12, :2002:12, :2004:12, :2007:9
      Register_inst134 <= _T_137[_T_2 == 8'h86 & write_0_en];	// <stdin>:2015:12, :2016:12, :2017:12, :2019:12, :2022:9
      Register_inst135 <= _T_138[_T_2 == 8'h87 & write_0_en];	// <stdin>:2030:12, :2031:12, :2032:12, :2034:12, :2037:9
      Register_inst136 <= _T_139[_T_2 == 8'h88 & write_0_en];	// <stdin>:2045:12, :2046:12, :2047:12, :2049:12, :2052:9
      Register_inst137 <= _T_140[_T_2 == 8'h89 & write_0_en];	// <stdin>:2060:12, :2061:12, :2062:12, :2064:12, :2067:9
      Register_inst138 <= _T_141[_T_2 == 8'h8A & write_0_en];	// <stdin>:2075:12, :2076:12, :2077:12, :2079:12, :2082:9
      Register_inst139 <= _T_142[_T_2 == 8'h8B & write_0_en];	// <stdin>:2090:12, :2091:12, :2092:12, :2094:12, :2097:9
      Register_inst140 <= _T_143[_T_2 == 8'h8C & write_0_en];	// <stdin>:2105:12, :2106:12, :2107:12, :2109:12, :2112:9
      Register_inst141 <= _T_144[_T_2 == 8'h8D & write_0_en];	// <stdin>:2120:12, :2121:12, :2122:12, :2124:12, :2127:9
      Register_inst142 <= _T_145[_T_2 == 8'h8E & write_0_en];	// <stdin>:2135:12, :2136:12, :2137:12, :2139:13, :2142:9
      Register_inst143 <= _T_146[_T_2 == 8'h8F & write_0_en];	// <stdin>:2150:13, :2151:13, :2152:13, :2154:13, :2157:9
      Register_inst144 <= _T_147[_T_2 == 8'h90 & write_0_en];	// <stdin>:2165:13, :2166:13, :2167:13, :2169:13, :2172:9
      Register_inst145 <= _T_148[_T_2 == 8'h91 & write_0_en];	// <stdin>:2180:13, :2181:13, :2182:13, :2184:13, :2187:9
      Register_inst146 <= _T_149[_T_2 == 8'h92 & write_0_en];	// <stdin>:2195:13, :2196:13, :2197:13, :2199:13, :2202:9
      Register_inst147 <= _T_150[_T_2 == 8'h93 & write_0_en];	// <stdin>:2210:13, :2211:13, :2212:13, :2214:13, :2217:9
      Register_inst148 <= _T_151[_T_2 == 8'h94 & write_0_en];	// <stdin>:2225:13, :2226:13, :2227:13, :2229:13, :2232:9
      Register_inst149 <= _T_152[_T_2 == 8'h95 & write_0_en];	// <stdin>:2240:13, :2241:13, :2242:13, :2244:13, :2247:9
      Register_inst150 <= _T_153[_T_2 == 8'h96 & write_0_en];	// <stdin>:2255:13, :2256:13, :2257:13, :2259:13, :2262:9
      Register_inst151 <= _T_154[_T_2 == 8'h97 & write_0_en];	// <stdin>:2270:13, :2271:13, :2272:13, :2274:13, :2277:9
      Register_inst152 <= _T_155[_T_2 == 8'h98 & write_0_en];	// <stdin>:2285:13, :2286:13, :2287:13, :2289:13, :2292:9
      Register_inst153 <= _T_156[_T_2 == 8'h99 & write_0_en];	// <stdin>:2300:13, :2301:13, :2302:13, :2304:13, :2307:9
      Register_inst154 <= _T_157[_T_2 == 8'h9A & write_0_en];	// <stdin>:2315:13, :2316:13, :2317:13, :2319:13, :2322:9
      Register_inst155 <= _T_158[_T_2 == 8'h9B & write_0_en];	// <stdin>:2330:13, :2331:13, :2332:13, :2334:13, :2337:9
      Register_inst156 <= _T_159[_T_2 == 8'h9C & write_0_en];	// <stdin>:2345:13, :2346:13, :2347:13, :2349:13, :2352:9
      Register_inst157 <= _T_160[_T_2 == 8'h9D & write_0_en];	// <stdin>:2360:13, :2361:13, :2362:13, :2364:13, :2367:9
      Register_inst158 <= _T_161[_T_2 == 8'h9E & write_0_en];	// <stdin>:2375:13, :2376:13, :2377:13, :2379:13, :2382:9
      Register_inst159 <= _T_162[_T_2 == 8'h9F & write_0_en];	// <stdin>:2390:13, :2391:13, :2392:13, :2394:13, :2397:9
      Register_inst160 <= _T_163[_T_2 == 8'hA0 & write_0_en];	// <stdin>:2405:13, :2406:13, :2407:13, :2409:13, :2412:9
      Register_inst161 <= _T_164[_T_2 == 8'hA1 & write_0_en];	// <stdin>:2420:13, :2421:13, :2422:13, :2424:13, :2427:9
      Register_inst162 <= _T_165[_T_2 == 8'hA2 & write_0_en];	// <stdin>:2435:13, :2436:13, :2437:13, :2439:13, :2442:9
      Register_inst163 <= _T_166[_T_2 == 8'hA3 & write_0_en];	// <stdin>:2450:13, :2451:13, :2452:13, :2454:13, :2457:9
      Register_inst164 <= _T_167[_T_2 == 8'hA4 & write_0_en];	// <stdin>:2465:13, :2466:13, :2467:13, :2469:13, :2472:9
      Register_inst165 <= _T_168[_T_2 == 8'hA5 & write_0_en];	// <stdin>:2480:13, :2481:13, :2482:13, :2484:13, :2487:9
      Register_inst166 <= _T_169[_T_2 == 8'hA6 & write_0_en];	// <stdin>:2495:13, :2496:13, :2497:13, :2499:13, :2502:9
      Register_inst167 <= _T_170[_T_2 == 8'hA7 & write_0_en];	// <stdin>:2510:13, :2511:13, :2512:13, :2514:13, :2517:9
      Register_inst168 <= _T_171[_T_2 == 8'hA8 & write_0_en];	// <stdin>:2525:13, :2526:13, :2527:13, :2529:13, :2532:9
      Register_inst169 <= _T_172[_T_2 == 8'hA9 & write_0_en];	// <stdin>:2540:13, :2541:13, :2542:13, :2544:13, :2547:9
      Register_inst170 <= _T_173[_T_2 == 8'hAA & write_0_en];	// <stdin>:2555:13, :2556:13, :2557:13, :2559:13, :2562:9
      Register_inst171 <= _T_174[_T_2 == 8'hAB & write_0_en];	// <stdin>:2570:13, :2571:13, :2572:13, :2574:13, :2577:9
      Register_inst172 <= _T_175[_T_2 == 8'hAC & write_0_en];	// <stdin>:2585:13, :2586:13, :2587:13, :2589:13, :2592:9
      Register_inst173 <= _T_176[_T_2 == 8'hAD & write_0_en];	// <stdin>:2600:13, :2601:13, :2602:13, :2604:13, :2607:9
      Register_inst174 <= _T_177[_T_2 == 8'hAE & write_0_en];	// <stdin>:2615:13, :2616:13, :2617:13, :2619:13, :2622:9
      Register_inst175 <= _T_178[_T_2 == 8'hAF & write_0_en];	// <stdin>:2630:13, :2631:13, :2632:13, :2634:13, :2637:9
      Register_inst176 <= _T_179[_T_2 == 8'hB0 & write_0_en];	// <stdin>:2645:13, :2646:13, :2647:13, :2649:13, :2652:9
      Register_inst177 <= _T_180[_T_2 == 8'hB1 & write_0_en];	// <stdin>:2660:13, :2661:13, :2662:13, :2664:13, :2667:9
      Register_inst178 <= _T_181[_T_2 == 8'hB2 & write_0_en];	// <stdin>:2675:13, :2676:13, :2677:13, :2679:13, :2682:9
      Register_inst179 <= _T_182[_T_2 == 8'hB3 & write_0_en];	// <stdin>:2690:13, :2691:13, :2692:13, :2694:13, :2697:9
      Register_inst180 <= _T_183[_T_2 == 8'hB4 & write_0_en];	// <stdin>:2705:13, :2706:13, :2707:13, :2709:13, :2712:9
      Register_inst181 <= _T_184[_T_2 == 8'hB5 & write_0_en];	// <stdin>:2720:13, :2721:13, :2722:13, :2724:13, :2727:9
      Register_inst182 <= _T_185[_T_2 == 8'hB6 & write_0_en];	// <stdin>:2735:13, :2736:13, :2737:13, :2739:13, :2742:9
      Register_inst183 <= _T_186[_T_2 == 8'hB7 & write_0_en];	// <stdin>:2750:13, :2751:13, :2752:13, :2754:13, :2757:9
      Register_inst184 <= _T_187[_T_2 == 8'hB8 & write_0_en];	// <stdin>:2765:13, :2766:13, :2767:13, :2769:13, :2772:9
      Register_inst185 <= _T_188[_T_2 == 8'hB9 & write_0_en];	// <stdin>:2780:13, :2781:13, :2782:13, :2784:13, :2787:9
      Register_inst186 <= _T_189[_T_2 == 8'hBA & write_0_en];	// <stdin>:2795:13, :2796:13, :2797:13, :2799:13, :2802:9
      Register_inst187 <= _T_190[_T_2 == 8'hBB & write_0_en];	// <stdin>:2810:13, :2811:13, :2812:13, :2814:13, :2817:9
      Register_inst188 <= _T_191[_T_2 == 8'hBC & write_0_en];	// <stdin>:2825:13, :2826:13, :2827:13, :2829:13, :2832:9
      Register_inst189 <= _T_192[_T_2 == 8'hBD & write_0_en];	// <stdin>:2840:13, :2841:13, :2842:13, :2844:13, :2847:9
      Register_inst190 <= _T_193[_T_2 == 8'hBE & write_0_en];	// <stdin>:2855:13, :2856:13, :2857:13, :2859:13, :2862:9
      Register_inst191 <= _T_194[_T_2 == 8'hBF & write_0_en];	// <stdin>:2870:13, :2871:13, :2872:13, :2874:13, :2877:9
      Register_inst192 <= _T_195[_T_2 == 8'hC0 & write_0_en];	// <stdin>:2885:13, :2886:13, :2887:13, :2889:13, :2892:9
      Register_inst193 <= _T_196[_T_2 == 8'hC1 & write_0_en];	// <stdin>:2900:13, :2901:13, :2902:13, :2904:13, :2907:9
      Register_inst194 <= _T_197[_T_2 == 8'hC2 & write_0_en];	// <stdin>:2915:13, :2916:13, :2917:13, :2919:13, :2922:9
      Register_inst195 <= _T_198[_T_2 == 8'hC3 & write_0_en];	// <stdin>:2930:13, :2931:13, :2932:13, :2934:13, :2937:9
      Register_inst196 <= _T_199[_T_2 == 8'hC4 & write_0_en];	// <stdin>:2945:13, :2946:13, :2947:13, :2949:13, :2952:9
      Register_inst197 <= _T_200[_T_2 == 8'hC5 & write_0_en];	// <stdin>:2960:13, :2961:13, :2962:13, :2964:13, :2967:9
      Register_inst198 <= _T_201[_T_2 == 8'hC6 & write_0_en];	// <stdin>:2975:13, :2976:13, :2977:13, :2979:13, :2982:9
      Register_inst199 <= _T_202[_T_2 == 8'hC7 & write_0_en];	// <stdin>:2990:13, :2991:13, :2992:13, :2994:13, :2997:9
      Register_inst200 <= _T_203[_T_2 == 8'hC8 & write_0_en];	// <stdin>:3005:13, :3006:13, :3007:13, :3009:13, :3012:9
      Register_inst201 <= _T_204[_T_2 == 8'hC9 & write_0_en];	// <stdin>:3020:13, :3021:13, :3022:13, :3024:13, :3027:9
      Register_inst202 <= _T_205[_T_2 == 8'hCA & write_0_en];	// <stdin>:3035:13, :3036:13, :3037:13, :3039:13, :3042:9
      Register_inst203 <= _T_206[_T_2 == 8'hCB & write_0_en];	// <stdin>:3050:13, :3051:13, :3052:13, :3054:13, :3057:9
      Register_inst204 <= _T_207[_T_2 == 8'hCC & write_0_en];	// <stdin>:3065:13, :3066:13, :3067:13, :3069:13, :3072:9
      Register_inst205 <= _T_208[_T_2 == 8'hCD & write_0_en];	// <stdin>:3080:13, :3081:13, :3082:13, :3084:13, :3087:9
      Register_inst206 <= _T_209[_T_2 == 8'hCE & write_0_en];	// <stdin>:3095:13, :3096:13, :3097:13, :3099:13, :3102:9
      Register_inst207 <= _T_210[_T_2 == 8'hCF & write_0_en];	// <stdin>:3110:13, :3111:13, :3112:13, :3114:13, :3117:9
      Register_inst208 <= _T_211[_T_2 == 8'hD0 & write_0_en];	// <stdin>:3125:13, :3126:13, :3127:13, :3129:13, :3132:9
      Register_inst209 <= _T_212[_T_2 == 8'hD1 & write_0_en];	// <stdin>:3140:13, :3141:13, :3142:13, :3144:13, :3147:9
      Register_inst210 <= _T_213[_T_2 == 8'hD2 & write_0_en];	// <stdin>:3155:13, :3156:13, :3157:13, :3159:13, :3162:9
      Register_inst211 <= _T_214[_T_2 == 8'hD3 & write_0_en];	// <stdin>:3170:13, :3171:13, :3172:13, :3174:13, :3177:9
      Register_inst212 <= _T_215[_T_2 == 8'hD4 & write_0_en];	// <stdin>:3185:13, :3186:13, :3187:13, :3189:13, :3192:9
      Register_inst213 <= _T_216[_T_2 == 8'hD5 & write_0_en];	// <stdin>:3200:13, :3201:13, :3202:13, :3204:13, :3207:9
      Register_inst214 <= _T_217[_T_2 == 8'hD6 & write_0_en];	// <stdin>:3215:13, :3216:13, :3217:13, :3219:13, :3222:9
      Register_inst215 <= _T_218[_T_2 == 8'hD7 & write_0_en];	// <stdin>:3230:13, :3231:13, :3232:13, :3234:13, :3237:9
      Register_inst216 <= _T_219[_T_2 == 8'hD8 & write_0_en];	// <stdin>:3245:13, :3246:13, :3247:13, :3249:13, :3252:9
      Register_inst217 <= _T_220[_T_2 == 8'hD9 & write_0_en];	// <stdin>:3260:13, :3261:13, :3262:13, :3264:13, :3267:9
      Register_inst218 <= _T_221[_T_2 == 8'hDA & write_0_en];	// <stdin>:3275:13, :3276:13, :3277:13, :3279:13, :3282:9
      Register_inst219 <= _T_222[_T_2 == 8'hDB & write_0_en];	// <stdin>:3290:13, :3291:13, :3292:13, :3294:13, :3297:9
      Register_inst220 <= _T_223[_T_2 == 8'hDC & write_0_en];	// <stdin>:3305:13, :3306:13, :3307:13, :3309:13, :3312:9
      Register_inst221 <= _T_224[_T_2 == 8'hDD & write_0_en];	// <stdin>:3320:13, :3321:13, :3322:13, :3324:13, :3327:9
      Register_inst222 <= _T_225[_T_2 == 8'hDE & write_0_en];	// <stdin>:3335:13, :3336:13, :3337:13, :3339:13, :3342:9
      Register_inst223 <= _T_226[_T_2 == 8'hDF & write_0_en];	// <stdin>:3350:13, :3351:13, :3352:13, :3354:13, :3357:9
      Register_inst224 <= _T_227[_T_2 == 8'hE0 & write_0_en];	// <stdin>:3365:13, :3366:13, :3367:13, :3369:13, :3372:9
      Register_inst225 <= _T_228[_T_2 == 8'hE1 & write_0_en];	// <stdin>:3380:13, :3381:13, :3382:13, :3384:13, :3387:9
      Register_inst226 <= _T_229[_T_2 == 8'hE2 & write_0_en];	// <stdin>:3395:13, :3396:13, :3397:13, :3399:13, :3402:9
      Register_inst227 <= _T_230[_T_2 == 8'hE3 & write_0_en];	// <stdin>:3410:13, :3411:13, :3412:13, :3414:13, :3417:9
      Register_inst228 <= _T_231[_T_2 == 8'hE4 & write_0_en];	// <stdin>:3425:13, :3426:13, :3427:13, :3429:13, :3432:9
      Register_inst229 <= _T_232[_T_2 == 8'hE5 & write_0_en];	// <stdin>:3440:13, :3441:13, :3442:13, :3444:13, :3447:9
      Register_inst230 <= _T_233[_T_2 == 8'hE6 & write_0_en];	// <stdin>:3455:13, :3456:13, :3457:13, :3459:13, :3462:9
      Register_inst231 <= _T_234[_T_2 == 8'hE7 & write_0_en];	// <stdin>:3470:13, :3471:13, :3472:13, :3474:13, :3477:9
      Register_inst232 <= _T_235[_T_2 == 8'hE8 & write_0_en];	// <stdin>:3485:13, :3486:13, :3487:13, :3489:13, :3492:9
      Register_inst233 <= _T_236[_T_2 == 8'hE9 & write_0_en];	// <stdin>:3500:13, :3501:13, :3502:13, :3504:13, :3507:9
      Register_inst234 <= _T_237[_T_2 == 8'hEA & write_0_en];	// <stdin>:3515:13, :3516:13, :3517:13, :3519:13, :3522:9
      Register_inst235 <= _T_238[_T_2 == 8'hEB & write_0_en];	// <stdin>:3530:13, :3531:13, :3532:13, :3534:13, :3537:9
      Register_inst236 <= _T_239[_T_2 == 8'hEC & write_0_en];	// <stdin>:3545:13, :3546:13, :3547:13, :3549:13, :3552:9
      Register_inst237 <= _T_240[_T_2 == 8'hED & write_0_en];	// <stdin>:3560:13, :3561:13, :3562:13, :3564:13, :3567:9
      Register_inst238 <= _T_241[_T_2 == 8'hEE & write_0_en];	// <stdin>:3575:13, :3576:13, :3577:13, :3579:13, :3582:9
      Register_inst239 <= _T_242[_T_2 == 8'hEF & write_0_en];	// <stdin>:3590:13, :3591:13, :3592:13, :3594:13, :3597:9
      Register_inst240 <= _T_243[_T_2 == 8'hF0 & write_0_en];	// <stdin>:3605:13, :3606:13, :3607:13, :3609:13, :3612:9
      Register_inst241 <= _T_244[_T_2 == 8'hF1 & write_0_en];	// <stdin>:3620:13, :3621:13, :3622:13, :3624:13, :3627:9
      Register_inst242 <= _T_245[_T_2 == 8'hF2 & write_0_en];	// <stdin>:3635:13, :3636:13, :3637:13, :3639:13, :3642:9
      Register_inst243 <= _T_246[_T_2 == 8'hF3 & write_0_en];	// <stdin>:3650:13, :3651:13, :3652:13, :3654:13, :3657:9
      Register_inst244 <= _T_247[_T_2 == 8'hF4 & write_0_en];	// <stdin>:3665:13, :3666:13, :3667:13, :3669:13, :3672:9
      Register_inst245 <= _T_248[_T_2 == 8'hF5 & write_0_en];	// <stdin>:3680:13, :3681:13, :3682:13, :3684:13, :3687:9
      Register_inst246 <= _T_249[_T_2 == 8'hF6 & write_0_en];	// <stdin>:3695:13, :3696:13, :3697:13, :3699:13, :3702:9
      Register_inst247 <= _T_250[_T_2 == 8'hF7 & write_0_en];	// <stdin>:3710:13, :3711:13, :3712:13, :3714:13, :3717:9
      Register_inst248 <= _T_251[_T_2 == 8'hF8 & write_0_en];	// <stdin>:3725:13, :3726:13, :3727:13, :3729:13, :3732:9
      Register_inst249 <= _T_252[_T_2 == 8'hF9 & write_0_en];	// <stdin>:3740:13, :3741:13, :3742:13, :3744:13, :3747:9
      Register_inst250 <= _T_253[_T_2 == 8'hFA & write_0_en];	// <stdin>:3755:13, :3756:13, :3757:13, :3759:13, :3762:9
      Register_inst251 <= _T_254[_T_2 == 8'hFB & write_0_en];	// <stdin>:3770:13, :3771:13, :3772:13, :3774:13, :3777:9
      Register_inst252 <= _T_255[_T_2 == 8'hFC & write_0_en];	// <stdin>:3785:13, :3786:13, :3787:13, :3789:13, :3792:9
      Register_inst253 <= _T_256[_T_2 == 8'hFD & write_0_en];	// <stdin>:3800:13, :3801:13, :3802:13, :3804:13, :3807:9
      Register_inst254 <= _T_257[_T_2 == 8'hFE & write_0_en];	// <stdin>:3815:13, :3816:13, :3817:13, :3819:13, :3822:9
      Register_inst255 <= _T_258[&_T_2 & write_0_en];	// <stdin>:3831:13, :3832:13, :3834:13, :3837:9
    end
  end // always_ff @(posedge or posedge)
  initial begin	// <stdin>:3841:5
    Register_inst0 = 32'h0;	// <stdin>:15:10, :17:9
    Register_inst1 = 32'h0;	// <stdin>:15:10, :32:9
    Register_inst2 = 32'h0;	// <stdin>:15:10, :47:9
    Register_inst3 = 32'h0;	// <stdin>:15:10, :62:9
    Register_inst4 = 32'h0;	// <stdin>:15:10, :77:9
    Register_inst5 = 32'h0;	// <stdin>:15:10, :92:9
    Register_inst6 = 32'h0;	// <stdin>:15:10, :107:9
    Register_inst7 = 32'h0;	// <stdin>:15:10, :122:9
    Register_inst8 = 32'h0;	// <stdin>:15:10, :137:9
    Register_inst9 = 32'h0;	// <stdin>:15:10, :152:9
    Register_inst10 = 32'h0;	// <stdin>:15:10, :167:9
    Register_inst11 = 32'h0;	// <stdin>:15:10, :182:9
    Register_inst12 = 32'h0;	// <stdin>:15:10, :197:9
    Register_inst13 = 32'h0;	// <stdin>:15:10, :212:9
    Register_inst14 = 32'h0;	// <stdin>:15:10, :227:9
    Register_inst15 = 32'h0;	// <stdin>:15:10, :242:9
    Register_inst16 = 32'h0;	// <stdin>:15:10, :257:9
    Register_inst17 = 32'h0;	// <stdin>:15:10, :272:9
    Register_inst18 = 32'h0;	// <stdin>:15:10, :287:9
    Register_inst19 = 32'h0;	// <stdin>:15:10, :302:9
    Register_inst20 = 32'h0;	// <stdin>:15:10, :317:9
    Register_inst21 = 32'h0;	// <stdin>:15:10, :332:9
    Register_inst22 = 32'h0;	// <stdin>:15:10, :347:9
    Register_inst23 = 32'h0;	// <stdin>:15:10, :362:9
    Register_inst24 = 32'h0;	// <stdin>:15:10, :377:9
    Register_inst25 = 32'h0;	// <stdin>:15:10, :392:9
    Register_inst26 = 32'h0;	// <stdin>:15:10, :407:9
    Register_inst27 = 32'h0;	// <stdin>:15:10, :422:9
    Register_inst28 = 32'h0;	// <stdin>:15:10, :437:9
    Register_inst29 = 32'h0;	// <stdin>:15:10, :452:9
    Register_inst30 = 32'h0;	// <stdin>:15:10, :467:9
    Register_inst31 = 32'h0;	// <stdin>:15:10, :482:9
    Register_inst32 = 32'h0;	// <stdin>:15:10, :497:9
    Register_inst33 = 32'h0;	// <stdin>:15:10, :512:9
    Register_inst34 = 32'h0;	// <stdin>:15:10, :527:9
    Register_inst35 = 32'h0;	// <stdin>:15:10, :542:9
    Register_inst36 = 32'h0;	// <stdin>:15:10, :557:9
    Register_inst37 = 32'h0;	// <stdin>:15:10, :572:9
    Register_inst38 = 32'h0;	// <stdin>:15:10, :587:9
    Register_inst39 = 32'h0;	// <stdin>:15:10, :602:9
    Register_inst40 = 32'h0;	// <stdin>:15:10, :617:9
    Register_inst41 = 32'h0;	// <stdin>:15:10, :632:9
    Register_inst42 = 32'h0;	// <stdin>:15:10, :647:9
    Register_inst43 = 32'h0;	// <stdin>:15:10, :662:9
    Register_inst44 = 32'h0;	// <stdin>:15:10, :677:9
    Register_inst45 = 32'h0;	// <stdin>:15:10, :692:9
    Register_inst46 = 32'h0;	// <stdin>:15:10, :707:9
    Register_inst47 = 32'h0;	// <stdin>:15:10, :722:9
    Register_inst48 = 32'h0;	// <stdin>:15:10, :737:9
    Register_inst49 = 32'h0;	// <stdin>:15:10, :752:9
    Register_inst50 = 32'h0;	// <stdin>:15:10, :767:9
    Register_inst51 = 32'h0;	// <stdin>:15:10, :782:9
    Register_inst52 = 32'h0;	// <stdin>:15:10, :797:9
    Register_inst53 = 32'h0;	// <stdin>:15:10, :812:9
    Register_inst54 = 32'h0;	// <stdin>:15:10, :827:9
    Register_inst55 = 32'h0;	// <stdin>:15:10, :842:9
    Register_inst56 = 32'h0;	// <stdin>:15:10, :857:9
    Register_inst57 = 32'h0;	// <stdin>:15:10, :872:9
    Register_inst58 = 32'h0;	// <stdin>:15:10, :887:9
    Register_inst59 = 32'h0;	// <stdin>:15:10, :902:9
    Register_inst60 = 32'h0;	// <stdin>:15:10, :917:9
    Register_inst61 = 32'h0;	// <stdin>:15:10, :932:9
    Register_inst62 = 32'h0;	// <stdin>:15:10, :947:9
    Register_inst63 = 32'h0;	// <stdin>:15:10, :962:9
    Register_inst64 = 32'h0;	// <stdin>:15:10, :977:9
    Register_inst65 = 32'h0;	// <stdin>:15:10, :992:9
    Register_inst66 = 32'h0;	// <stdin>:15:10, :1007:9
    Register_inst67 = 32'h0;	// <stdin>:15:10, :1022:9
    Register_inst68 = 32'h0;	// <stdin>:15:10, :1037:9
    Register_inst69 = 32'h0;	// <stdin>:15:10, :1052:9
    Register_inst70 = 32'h0;	// <stdin>:15:10, :1067:9
    Register_inst71 = 32'h0;	// <stdin>:15:10, :1082:9
    Register_inst72 = 32'h0;	// <stdin>:15:10, :1097:9
    Register_inst73 = 32'h0;	// <stdin>:15:10, :1112:9
    Register_inst74 = 32'h0;	// <stdin>:15:10, :1127:9
    Register_inst75 = 32'h0;	// <stdin>:15:10, :1142:9
    Register_inst76 = 32'h0;	// <stdin>:15:10, :1157:9
    Register_inst77 = 32'h0;	// <stdin>:15:10, :1172:9
    Register_inst78 = 32'h0;	// <stdin>:15:10, :1187:9
    Register_inst79 = 32'h0;	// <stdin>:15:10, :1202:9
    Register_inst80 = 32'h0;	// <stdin>:15:10, :1217:9
    Register_inst81 = 32'h0;	// <stdin>:15:10, :1232:9
    Register_inst82 = 32'h0;	// <stdin>:15:10, :1247:9
    Register_inst83 = 32'h0;	// <stdin>:15:10, :1262:9
    Register_inst84 = 32'h0;	// <stdin>:15:10, :1277:9
    Register_inst85 = 32'h0;	// <stdin>:15:10, :1292:9
    Register_inst86 = 32'h0;	// <stdin>:15:10, :1307:9
    Register_inst87 = 32'h0;	// <stdin>:15:10, :1322:9
    Register_inst88 = 32'h0;	// <stdin>:15:10, :1337:9
    Register_inst89 = 32'h0;	// <stdin>:15:10, :1352:9
    Register_inst90 = 32'h0;	// <stdin>:15:10, :1367:9
    Register_inst91 = 32'h0;	// <stdin>:15:10, :1382:9
    Register_inst92 = 32'h0;	// <stdin>:15:10, :1397:9
    Register_inst93 = 32'h0;	// <stdin>:15:10, :1412:9
    Register_inst94 = 32'h0;	// <stdin>:15:10, :1427:9
    Register_inst95 = 32'h0;	// <stdin>:15:10, :1442:9
    Register_inst96 = 32'h0;	// <stdin>:15:10, :1457:9
    Register_inst97 = 32'h0;	// <stdin>:15:10, :1472:9
    Register_inst98 = 32'h0;	// <stdin>:15:10, :1487:9
    Register_inst99 = 32'h0;	// <stdin>:15:10, :1502:9
    Register_inst100 = 32'h0;	// <stdin>:15:10, :1517:9
    Register_inst101 = 32'h0;	// <stdin>:15:10, :1532:9
    Register_inst102 = 32'h0;	// <stdin>:15:10, :1547:9
    Register_inst103 = 32'h0;	// <stdin>:15:10, :1562:9
    Register_inst104 = 32'h0;	// <stdin>:15:10, :1577:9
    Register_inst105 = 32'h0;	// <stdin>:15:10, :1592:9
    Register_inst106 = 32'h0;	// <stdin>:15:10, :1607:9
    Register_inst107 = 32'h0;	// <stdin>:15:10, :1622:9
    Register_inst108 = 32'h0;	// <stdin>:15:10, :1637:9
    Register_inst109 = 32'h0;	// <stdin>:15:10, :1652:9
    Register_inst110 = 32'h0;	// <stdin>:15:10, :1667:9
    Register_inst111 = 32'h0;	// <stdin>:15:10, :1682:9
    Register_inst112 = 32'h0;	// <stdin>:15:10, :1697:9
    Register_inst113 = 32'h0;	// <stdin>:15:10, :1712:9
    Register_inst114 = 32'h0;	// <stdin>:15:10, :1727:9
    Register_inst115 = 32'h0;	// <stdin>:15:10, :1742:9
    Register_inst116 = 32'h0;	// <stdin>:15:10, :1757:9
    Register_inst117 = 32'h0;	// <stdin>:15:10, :1772:9
    Register_inst118 = 32'h0;	// <stdin>:15:10, :1787:9
    Register_inst119 = 32'h0;	// <stdin>:15:10, :1802:9
    Register_inst120 = 32'h0;	// <stdin>:15:10, :1817:9
    Register_inst121 = 32'h0;	// <stdin>:15:10, :1832:9
    Register_inst122 = 32'h0;	// <stdin>:15:10, :1847:9
    Register_inst123 = 32'h0;	// <stdin>:15:10, :1862:9
    Register_inst124 = 32'h0;	// <stdin>:15:10, :1877:9
    Register_inst125 = 32'h0;	// <stdin>:15:10, :1892:9
    Register_inst126 = 32'h0;	// <stdin>:15:10, :1907:9
    Register_inst127 = 32'h0;	// <stdin>:15:10, :1922:9
    Register_inst128 = 32'h0;	// <stdin>:15:10, :1937:9
    Register_inst129 = 32'h0;	// <stdin>:15:10, :1952:9
    Register_inst130 = 32'h0;	// <stdin>:15:10, :1967:9
    Register_inst131 = 32'h0;	// <stdin>:15:10, :1982:9
    Register_inst132 = 32'h0;	// <stdin>:15:10, :1997:9
    Register_inst133 = 32'h0;	// <stdin>:15:10, :2012:9
    Register_inst134 = 32'h0;	// <stdin>:15:10, :2027:9
    Register_inst135 = 32'h0;	// <stdin>:15:10, :2042:9
    Register_inst136 = 32'h0;	// <stdin>:15:10, :2057:9
    Register_inst137 = 32'h0;	// <stdin>:15:10, :2072:9
    Register_inst138 = 32'h0;	// <stdin>:15:10, :2087:9
    Register_inst139 = 32'h0;	// <stdin>:15:10, :2102:9
    Register_inst140 = 32'h0;	// <stdin>:15:10, :2117:9
    Register_inst141 = 32'h0;	// <stdin>:15:10, :2132:9
    Register_inst142 = 32'h0;	// <stdin>:15:10, :2147:9
    Register_inst143 = 32'h0;	// <stdin>:15:10, :2162:9
    Register_inst144 = 32'h0;	// <stdin>:15:10, :2177:9
    Register_inst145 = 32'h0;	// <stdin>:15:10, :2192:9
    Register_inst146 = 32'h0;	// <stdin>:15:10, :2207:9
    Register_inst147 = 32'h0;	// <stdin>:15:10, :2222:9
    Register_inst148 = 32'h0;	// <stdin>:15:10, :2237:9
    Register_inst149 = 32'h0;	// <stdin>:15:10, :2252:9
    Register_inst150 = 32'h0;	// <stdin>:15:10, :2267:9
    Register_inst151 = 32'h0;	// <stdin>:15:10, :2282:9
    Register_inst152 = 32'h0;	// <stdin>:15:10, :2297:9
    Register_inst153 = 32'h0;	// <stdin>:15:10, :2312:9
    Register_inst154 = 32'h0;	// <stdin>:15:10, :2327:9
    Register_inst155 = 32'h0;	// <stdin>:15:10, :2342:9
    Register_inst156 = 32'h0;	// <stdin>:15:10, :2357:9
    Register_inst157 = 32'h0;	// <stdin>:15:10, :2372:9
    Register_inst158 = 32'h0;	// <stdin>:15:10, :2387:9
    Register_inst159 = 32'h0;	// <stdin>:15:10, :2402:9
    Register_inst160 = 32'h0;	// <stdin>:15:10, :2417:9
    Register_inst161 = 32'h0;	// <stdin>:15:10, :2432:9
    Register_inst162 = 32'h0;	// <stdin>:15:10, :2447:9
    Register_inst163 = 32'h0;	// <stdin>:15:10, :2462:9
    Register_inst164 = 32'h0;	// <stdin>:15:10, :2477:9
    Register_inst165 = 32'h0;	// <stdin>:15:10, :2492:9
    Register_inst166 = 32'h0;	// <stdin>:15:10, :2507:9
    Register_inst167 = 32'h0;	// <stdin>:15:10, :2522:9
    Register_inst168 = 32'h0;	// <stdin>:15:10, :2537:9
    Register_inst169 = 32'h0;	// <stdin>:15:10, :2552:9
    Register_inst170 = 32'h0;	// <stdin>:15:10, :2567:9
    Register_inst171 = 32'h0;	// <stdin>:15:10, :2582:9
    Register_inst172 = 32'h0;	// <stdin>:15:10, :2597:9
    Register_inst173 = 32'h0;	// <stdin>:15:10, :2612:9
    Register_inst174 = 32'h0;	// <stdin>:15:10, :2627:9
    Register_inst175 = 32'h0;	// <stdin>:15:10, :2642:9
    Register_inst176 = 32'h0;	// <stdin>:15:10, :2657:9
    Register_inst177 = 32'h0;	// <stdin>:15:10, :2672:9
    Register_inst178 = 32'h0;	// <stdin>:15:10, :2687:9
    Register_inst179 = 32'h0;	// <stdin>:15:10, :2702:9
    Register_inst180 = 32'h0;	// <stdin>:15:10, :2717:9
    Register_inst181 = 32'h0;	// <stdin>:15:10, :2732:9
    Register_inst182 = 32'h0;	// <stdin>:15:10, :2747:9
    Register_inst183 = 32'h0;	// <stdin>:15:10, :2762:9
    Register_inst184 = 32'h0;	// <stdin>:15:10, :2777:9
    Register_inst185 = 32'h0;	// <stdin>:15:10, :2792:9
    Register_inst186 = 32'h0;	// <stdin>:15:10, :2807:9
    Register_inst187 = 32'h0;	// <stdin>:15:10, :2822:9
    Register_inst188 = 32'h0;	// <stdin>:15:10, :2837:9
    Register_inst189 = 32'h0;	// <stdin>:15:10, :2852:9
    Register_inst190 = 32'h0;	// <stdin>:15:10, :2867:9
    Register_inst191 = 32'h0;	// <stdin>:15:10, :2882:9
    Register_inst192 = 32'h0;	// <stdin>:15:10, :2897:9
    Register_inst193 = 32'h0;	// <stdin>:15:10, :2912:9
    Register_inst194 = 32'h0;	// <stdin>:15:10, :2927:9
    Register_inst195 = 32'h0;	// <stdin>:15:10, :2942:9
    Register_inst196 = 32'h0;	// <stdin>:15:10, :2957:9
    Register_inst197 = 32'h0;	// <stdin>:15:10, :2972:9
    Register_inst198 = 32'h0;	// <stdin>:15:10, :2987:9
    Register_inst199 = 32'h0;	// <stdin>:15:10, :3002:9
    Register_inst200 = 32'h0;	// <stdin>:15:10, :3017:9
    Register_inst201 = 32'h0;	// <stdin>:15:10, :3032:9
    Register_inst202 = 32'h0;	// <stdin>:15:10, :3047:9
    Register_inst203 = 32'h0;	// <stdin>:15:10, :3062:9
    Register_inst204 = 32'h0;	// <stdin>:15:10, :3077:9
    Register_inst205 = 32'h0;	// <stdin>:15:10, :3092:9
    Register_inst206 = 32'h0;	// <stdin>:15:10, :3107:9
    Register_inst207 = 32'h0;	// <stdin>:15:10, :3122:9
    Register_inst208 = 32'h0;	// <stdin>:15:10, :3137:9
    Register_inst209 = 32'h0;	// <stdin>:15:10, :3152:9
    Register_inst210 = 32'h0;	// <stdin>:15:10, :3167:9
    Register_inst211 = 32'h0;	// <stdin>:15:10, :3182:9
    Register_inst212 = 32'h0;	// <stdin>:15:10, :3197:9
    Register_inst213 = 32'h0;	// <stdin>:15:10, :3212:9
    Register_inst214 = 32'h0;	// <stdin>:15:10, :3227:9
    Register_inst215 = 32'h0;	// <stdin>:15:10, :3242:9
    Register_inst216 = 32'h0;	// <stdin>:15:10, :3257:9
    Register_inst217 = 32'h0;	// <stdin>:15:10, :3272:9
    Register_inst218 = 32'h0;	// <stdin>:15:10, :3287:9
    Register_inst219 = 32'h0;	// <stdin>:15:10, :3302:9
    Register_inst220 = 32'h0;	// <stdin>:15:10, :3317:9
    Register_inst221 = 32'h0;	// <stdin>:15:10, :3332:9
    Register_inst222 = 32'h0;	// <stdin>:15:10, :3347:9
    Register_inst223 = 32'h0;	// <stdin>:15:10, :3362:9
    Register_inst224 = 32'h0;	// <stdin>:15:10, :3377:9
    Register_inst225 = 32'h0;	// <stdin>:15:10, :3392:9
    Register_inst226 = 32'h0;	// <stdin>:15:10, :3407:9
    Register_inst227 = 32'h0;	// <stdin>:15:10, :3422:9
    Register_inst228 = 32'h0;	// <stdin>:15:10, :3437:9
    Register_inst229 = 32'h0;	// <stdin>:15:10, :3452:9
    Register_inst230 = 32'h0;	// <stdin>:15:10, :3467:9
    Register_inst231 = 32'h0;	// <stdin>:15:10, :3482:9
    Register_inst232 = 32'h0;	// <stdin>:15:10, :3497:9
    Register_inst233 = 32'h0;	// <stdin>:15:10, :3512:9
    Register_inst234 = 32'h0;	// <stdin>:15:10, :3527:9
    Register_inst235 = 32'h0;	// <stdin>:15:10, :3542:9
    Register_inst236 = 32'h0;	// <stdin>:15:10, :3557:9
    Register_inst237 = 32'h0;	// <stdin>:15:10, :3572:9
    Register_inst238 = 32'h0;	// <stdin>:15:10, :3587:9
    Register_inst239 = 32'h0;	// <stdin>:15:10, :3602:9
    Register_inst240 = 32'h0;	// <stdin>:15:10, :3617:9
    Register_inst241 = 32'h0;	// <stdin>:15:10, :3632:9
    Register_inst242 = 32'h0;	// <stdin>:15:10, :3647:9
    Register_inst243 = 32'h0;	// <stdin>:15:10, :3662:9
    Register_inst244 = 32'h0;	// <stdin>:15:10, :3677:9
    Register_inst245 = 32'h0;	// <stdin>:15:10, :3692:9
    Register_inst246 = 32'h0;	// <stdin>:15:10, :3707:9
    Register_inst247 = 32'h0;	// <stdin>:15:10, :3722:9
    Register_inst248 = 32'h0;	// <stdin>:15:10, :3737:9
    Register_inst249 = 32'h0;	// <stdin>:15:10, :3752:9
    Register_inst250 = 32'h0;	// <stdin>:15:10, :3767:9
    Register_inst251 = 32'h0;	// <stdin>:15:10, :3782:9
    Register_inst252 = 32'h0;	// <stdin>:15:10, :3797:9
    Register_inst253 = 32'h0;	// <stdin>:15:10, :3812:9
    Register_inst254 = 32'h0;	// <stdin>:15:10, :3827:9
    Register_inst255 = 32'h0;	// <stdin>:15:10, :3842:9
  end // initial
  wire [255:0][31:0] _T = {{Register_inst0}, {Register_inst1}, {Register_inst2}, {Register_inst3}, {Register_inst4},
                {Register_inst5}, {Register_inst6}, {Register_inst7}, {Register_inst8}, {Register_inst9},
                {Register_inst10}, {Register_inst11}, {Register_inst12}, {Register_inst13},
                {Register_inst14}, {Register_inst15}, {Register_inst16}, {Register_inst17},
                {Register_inst18}, {Register_inst19}, {Register_inst20}, {Register_inst21},
                {Register_inst22}, {Register_inst23}, {Register_inst24}, {Register_inst25},
                {Register_inst26}, {Register_inst27}, {Register_inst28}, {Register_inst29},
                {Register_inst30}, {Register_inst31}, {Register_inst32}, {Register_inst33},
                {Register_inst34}, {Register_inst35}, {Register_inst36}, {Register_inst37},
                {Register_inst38}, {Register_inst39}, {Register_inst40}, {Register_inst41},
                {Register_inst42}, {Register_inst43}, {Register_inst44}, {Register_inst45},
                {Register_inst46}, {Register_inst47}, {Register_inst48}, {Register_inst49},
                {Register_inst50}, {Register_inst51}, {Register_inst52}, {Register_inst53},
                {Register_inst54}, {Register_inst55}, {Register_inst56}, {Register_inst57},
                {Register_inst58}, {Register_inst59}, {Register_inst60}, {Register_inst61},
                {Register_inst62}, {Register_inst63}, {Register_inst64}, {Register_inst65},
                {Register_inst66}, {Register_inst67}, {Register_inst68}, {Register_inst69},
                {Register_inst70}, {Register_inst71}, {Register_inst72}, {Register_inst73},
                {Register_inst74}, {Register_inst75}, {Register_inst76}, {Register_inst77},
                {Register_inst78}, {Register_inst79}, {Register_inst80}, {Register_inst81},
                {Register_inst82}, {Register_inst83}, {Register_inst84}, {Register_inst85},
                {Register_inst86}, {Register_inst87}, {Register_inst88}, {Register_inst89},
                {Register_inst90}, {Register_inst91}, {Register_inst92}, {Register_inst93},
                {Register_inst94}, {Register_inst95}, {Register_inst96}, {Register_inst97},
                {Register_inst98}, {Register_inst99}, {Register_inst100}, {Register_inst101},
                {Register_inst102}, {Register_inst103}, {Register_inst104}, {Register_inst105},
                {Register_inst106}, {Register_inst107}, {Register_inst108}, {Register_inst109},
                {Register_inst110}, {Register_inst111}, {Register_inst112}, {Register_inst113},
                {Register_inst114}, {Register_inst115}, {Register_inst116}, {Register_inst117},
                {Register_inst118}, {Register_inst119}, {Register_inst120}, {Register_inst121},
                {Register_inst122}, {Register_inst123}, {Register_inst124}, {Register_inst125},
                {Register_inst126}, {Register_inst127}, {Register_inst128}, {Register_inst129},
                {Register_inst130}, {Register_inst131}, {Register_inst132}, {Register_inst133},
                {Register_inst134}, {Register_inst135}, {Register_inst136}, {Register_inst137},
                {Register_inst138}, {Register_inst139}, {Register_inst140}, {Register_inst141},
                {Register_inst142}, {Register_inst143}, {Register_inst144}, {Register_inst145},
                {Register_inst146}, {Register_inst147}, {Register_inst148}, {Register_inst149},
                {Register_inst150}, {Register_inst151}, {Register_inst152}, {Register_inst153},
                {Register_inst154}, {Register_inst155}, {Register_inst156}, {Register_inst157},
                {Register_inst158}, {Register_inst159}, {Register_inst160}, {Register_inst161},
                {Register_inst162}, {Register_inst163}, {Register_inst164}, {Register_inst165},
                {Register_inst166}, {Register_inst167}, {Register_inst168}, {Register_inst169},
                {Register_inst170}, {Register_inst171}, {Register_inst172}, {Register_inst173},
                {Register_inst174}, {Register_inst175}, {Register_inst176}, {Register_inst177},
                {Register_inst178}, {Register_inst179}, {Register_inst180}, {Register_inst181},
                {Register_inst182}, {Register_inst183}, {Register_inst184}, {Register_inst185},
                {Register_inst186}, {Register_inst187}, {Register_inst188}, {Register_inst189},
                {Register_inst190}, {Register_inst191}, {Register_inst192}, {Register_inst193},
                {Register_inst194}, {Register_inst195}, {Register_inst196}, {Register_inst197},
                {Register_inst198}, {Register_inst199}, {Register_inst200}, {Register_inst201},
                {Register_inst202}, {Register_inst203}, {Register_inst204}, {Register_inst205},
                {Register_inst206}, {Register_inst207}, {Register_inst208}, {Register_inst209},
                {Register_inst210}, {Register_inst211}, {Register_inst212}, {Register_inst213},
                {Register_inst214}, {Register_inst215}, {Register_inst216}, {Register_inst217},
                {Register_inst218}, {Register_inst219}, {Register_inst220}, {Register_inst221},
                {Register_inst222}, {Register_inst223}, {Register_inst224}, {Register_inst225},
                {Register_inst226}, {Register_inst227}, {Register_inst228}, {Register_inst229},
                {Register_inst230}, {Register_inst231}, {Register_inst232}, {Register_inst233},
                {Register_inst234}, {Register_inst235}, {Register_inst236}, {Register_inst237},
                {Register_inst238}, {Register_inst239}, {Register_inst240}, {Register_inst241},
                {Register_inst242}, {Register_inst243}, {Register_inst244}, {Register_inst245},
                {Register_inst246}, {Register_inst247}, {Register_inst248}, {Register_inst249},
                {Register_inst250}, {Register_inst251}, {Register_inst252}, {Register_inst253},
                {Register_inst254}, {Register_inst255}};	// <stdin>:19:10, :34:11, :49:11, :64:11, :79:11, :94:11, :109:11, :124:11, :139:11, :154:11, :169:11, :184:11, :199:11, :214:11, :229:12, :244:12, :259:12, :274:12, :289:12, :304:12, :319:12, :334:12, :349:12, :364:12, :379:12, :394:12, :409:12, :424:12, :439:12, :454:12, :469:12, :484:12, :499:12, :514:12, :529:12, :544:12, :559:12, :574:12, :589:12, :604:12, :619:12, :634:12, :649:12, :664:12, :679:12, :694:12, :709:12, :724:12, :739:12, :754:12, :769:12, :784:12, :799:12, :814:12, :829:12, :844:12, :859:12, :874:12, :889:12, :904:12, :919:12, :934:12, :949:12, :964:12, :979:12, :994:12, :1009:12, :1024:12, :1039:12, :1054:12, :1069:12, :1084:12, :1099:12, :1114:12, :1129:12, :1144:12, :1159:12, :1174:12, :1189:12, :1204:12, :1219:12, :1234:12, :1249:12, :1264:12, :1279:12, :1294:12, :1309:12, :1324:12, :1339:12, :1354:12, :1369:12, :1384:12, :1399:12, :1414:12, :1429:12, :1444:12, :1459:12, :1474:12, :1489:12, :1504:12, :1519:12, :1534:12, :1549:12, :1564:12, :1579:12, :1594:12, :1609:12, :1624:12, :1639:12, :1654:12, :1669:12, :1684:12, :1699:12, :1714:12, :1729:12, :1744:12, :1759:12, :1774:12, :1789:12, :1804:12, :1819:12, :1834:12, :1849:12, :1864:12, :1879:12, :1894:12, :1909:12, :1924:12, :1939:12, :1954:12, :1969:12, :1984:12, :1999:12, :2014:12, :2029:12, :2044:12, :2059:12, :2074:12, :2089:12, :2104:12, :2119:12, :2134:12, :2149:13, :2164:13, :2179:13, :2194:13, :2209:13, :2224:13, :2239:13, :2254:13, :2269:13, :2284:13, :2299:13, :2314:13, :2329:13, :2344:13, :2359:13, :2374:13, :2389:13, :2404:13, :2419:13, :2434:13, :2449:13, :2464:13, :2479:13, :2494:13, :2509:13, :2524:13, :2539:13, :2554:13, :2569:13, :2584:13, :2599:13, :2614:13, :2629:13, :2644:13, :2659:13, :2674:13, :2689:13, :2704:13, :2719:13, :2734:13, :2749:13, :2764:13, :2779:13, :2794:13, :2809:13, :2824:13, :2839:13, :2854:13, :2869:13, :2884:13, :2899:13, :2914:13, :2929:13, :2944:13, :2959:13, :2974:13, :2989:13, :3004:13, :3019:13, :3034:13, :3049:13, :3064:13, :3079:13, :3094:13, :3109:13, :3124:13, :3139:13, :3154:13, :3169:13, :3184:13, :3199:13, :3214:13, :3229:13, :3244:13, :3259:13, :3274:13, :3289:13, :3304:13, :3319:13, :3334:13, :3349:13, :3364:13, :3379:13, :3394:13, :3409:13, :3424:13, :3439:13, :3454:13, :3469:13, :3484:13, :3499:13, :3514:13, :3529:13, :3544:13, :3559:13, :3574:13, :3589:13, :3604:13, :3619:13, :3634:13, :3649:13, :3664:13, :3679:13, :3694:13, :3709:13, :3724:13, :3739:13, :3754:13, :3769:13, :3784:13, :3799:13, :3814:13, :3829:13, :3844:13, :3845:13
  wire [255:0][31:0] _T_0 = {{Register_inst0}, {Register_inst1}, {Register_inst2}, {Register_inst3}, {Register_inst4},
                {Register_inst5}, {Register_inst6}, {Register_inst7}, {Register_inst8}, {Register_inst9},
                {Register_inst10}, {Register_inst11}, {Register_inst12}, {Register_inst13},
                {Register_inst14}, {Register_inst15}, {Register_inst16}, {Register_inst17},
                {Register_inst18}, {Register_inst19}, {Register_inst20}, {Register_inst21},
                {Register_inst22}, {Register_inst23}, {Register_inst24}, {Register_inst25},
                {Register_inst26}, {Register_inst27}, {Register_inst28}, {Register_inst29},
                {Register_inst30}, {Register_inst31}, {Register_inst32}, {Register_inst33},
                {Register_inst34}, {Register_inst35}, {Register_inst36}, {Register_inst37},
                {Register_inst38}, {Register_inst39}, {Register_inst40}, {Register_inst41},
                {Register_inst42}, {Register_inst43}, {Register_inst44}, {Register_inst45},
                {Register_inst46}, {Register_inst47}, {Register_inst48}, {Register_inst49},
                {Register_inst50}, {Register_inst51}, {Register_inst52}, {Register_inst53},
                {Register_inst54}, {Register_inst55}, {Register_inst56}, {Register_inst57},
                {Register_inst58}, {Register_inst59}, {Register_inst60}, {Register_inst61},
                {Register_inst62}, {Register_inst63}, {Register_inst64}, {Register_inst65},
                {Register_inst66}, {Register_inst67}, {Register_inst68}, {Register_inst69},
                {Register_inst70}, {Register_inst71}, {Register_inst72}, {Register_inst73},
                {Register_inst74}, {Register_inst75}, {Register_inst76}, {Register_inst77},
                {Register_inst78}, {Register_inst79}, {Register_inst80}, {Register_inst81},
                {Register_inst82}, {Register_inst83}, {Register_inst84}, {Register_inst85},
                {Register_inst86}, {Register_inst87}, {Register_inst88}, {Register_inst89},
                {Register_inst90}, {Register_inst91}, {Register_inst92}, {Register_inst93},
                {Register_inst94}, {Register_inst95}, {Register_inst96}, {Register_inst97},
                {Register_inst98}, {Register_inst99}, {Register_inst100}, {Register_inst101},
                {Register_inst102}, {Register_inst103}, {Register_inst104}, {Register_inst105},
                {Register_inst106}, {Register_inst107}, {Register_inst108}, {Register_inst109},
                {Register_inst110}, {Register_inst111}, {Register_inst112}, {Register_inst113},
                {Register_inst114}, {Register_inst115}, {Register_inst116}, {Register_inst117},
                {Register_inst118}, {Register_inst119}, {Register_inst120}, {Register_inst121},
                {Register_inst122}, {Register_inst123}, {Register_inst124}, {Register_inst125},
                {Register_inst126}, {Register_inst127}, {Register_inst128}, {Register_inst129},
                {Register_inst130}, {Register_inst131}, {Register_inst132}, {Register_inst133},
                {Register_inst134}, {Register_inst135}, {Register_inst136}, {Register_inst137},
                {Register_inst138}, {Register_inst139}, {Register_inst140}, {Register_inst141},
                {Register_inst142}, {Register_inst143}, {Register_inst144}, {Register_inst145},
                {Register_inst146}, {Register_inst147}, {Register_inst148}, {Register_inst149},
                {Register_inst150}, {Register_inst151}, {Register_inst152}, {Register_inst153},
                {Register_inst154}, {Register_inst155}, {Register_inst156}, {Register_inst157},
                {Register_inst158}, {Register_inst159}, {Register_inst160}, {Register_inst161},
                {Register_inst162}, {Register_inst163}, {Register_inst164}, {Register_inst165},
                {Register_inst166}, {Register_inst167}, {Register_inst168}, {Register_inst169},
                {Register_inst170}, {Register_inst171}, {Register_inst172}, {Register_inst173},
                {Register_inst174}, {Register_inst175}, {Register_inst176}, {Register_inst177},
                {Register_inst178}, {Register_inst179}, {Register_inst180}, {Register_inst181},
                {Register_inst182}, {Register_inst183}, {Register_inst184}, {Register_inst185},
                {Register_inst186}, {Register_inst187}, {Register_inst188}, {Register_inst189},
                {Register_inst190}, {Register_inst191}, {Register_inst192}, {Register_inst193},
                {Register_inst194}, {Register_inst195}, {Register_inst196}, {Register_inst197},
                {Register_inst198}, {Register_inst199}, {Register_inst200}, {Register_inst201},
                {Register_inst202}, {Register_inst203}, {Register_inst204}, {Register_inst205},
                {Register_inst206}, {Register_inst207}, {Register_inst208}, {Register_inst209},
                {Register_inst210}, {Register_inst211}, {Register_inst212}, {Register_inst213},
                {Register_inst214}, {Register_inst215}, {Register_inst216}, {Register_inst217},
                {Register_inst218}, {Register_inst219}, {Register_inst220}, {Register_inst221},
                {Register_inst222}, {Register_inst223}, {Register_inst224}, {Register_inst225},
                {Register_inst226}, {Register_inst227}, {Register_inst228}, {Register_inst229},
                {Register_inst230}, {Register_inst231}, {Register_inst232}, {Register_inst233},
                {Register_inst234}, {Register_inst235}, {Register_inst236}, {Register_inst237},
                {Register_inst238}, {Register_inst239}, {Register_inst240}, {Register_inst241},
                {Register_inst242}, {Register_inst243}, {Register_inst244}, {Register_inst245},
                {Register_inst246}, {Register_inst247}, {Register_inst248}, {Register_inst249},
                {Register_inst250}, {Register_inst251}, {Register_inst252}, {Register_inst253},
                {Register_inst254}, {Register_inst255}};	// <stdin>:19:10, :34:11, :49:11, :64:11, :79:11, :94:11, :109:11, :124:11, :139:11, :154:11, :169:11, :184:11, :199:11, :214:11, :229:12, :244:12, :259:12, :274:12, :289:12, :304:12, :319:12, :334:12, :349:12, :364:12, :379:12, :394:12, :409:12, :424:12, :439:12, :454:12, :469:12, :484:12, :499:12, :514:12, :529:12, :544:12, :559:12, :574:12, :589:12, :604:12, :619:12, :634:12, :649:12, :664:12, :679:12, :694:12, :709:12, :724:12, :739:12, :754:12, :769:12, :784:12, :799:12, :814:12, :829:12, :844:12, :859:12, :874:12, :889:12, :904:12, :919:12, :934:12, :949:12, :964:12, :979:12, :994:12, :1009:12, :1024:12, :1039:12, :1054:12, :1069:12, :1084:12, :1099:12, :1114:12, :1129:12, :1144:12, :1159:12, :1174:12, :1189:12, :1204:12, :1219:12, :1234:12, :1249:12, :1264:12, :1279:12, :1294:12, :1309:12, :1324:12, :1339:12, :1354:12, :1369:12, :1384:12, :1399:12, :1414:12, :1429:12, :1444:12, :1459:12, :1474:12, :1489:12, :1504:12, :1519:12, :1534:12, :1549:12, :1564:12, :1579:12, :1594:12, :1609:12, :1624:12, :1639:12, :1654:12, :1669:12, :1684:12, :1699:12, :1714:12, :1729:12, :1744:12, :1759:12, :1774:12, :1789:12, :1804:12, :1819:12, :1834:12, :1849:12, :1864:12, :1879:12, :1894:12, :1909:12, :1924:12, :1939:12, :1954:12, :1969:12, :1984:12, :1999:12, :2014:12, :2029:12, :2044:12, :2059:12, :2074:12, :2089:12, :2104:12, :2119:12, :2134:12, :2149:13, :2164:13, :2179:13, :2194:13, :2209:13, :2224:13, :2239:13, :2254:13, :2269:13, :2284:13, :2299:13, :2314:13, :2329:13, :2344:13, :2359:13, :2374:13, :2389:13, :2404:13, :2419:13, :2434:13, :2449:13, :2464:13, :2479:13, :2494:13, :2509:13, :2524:13, :2539:13, :2554:13, :2569:13, :2584:13, :2599:13, :2614:13, :2629:13, :2644:13, :2659:13, :2674:13, :2689:13, :2704:13, :2719:13, :2734:13, :2749:13, :2764:13, :2779:13, :2794:13, :2809:13, :2824:13, :2839:13, :2854:13, :2869:13, :2884:13, :2899:13, :2914:13, :2929:13, :2944:13, :2959:13, :2974:13, :2989:13, :3004:13, :3019:13, :3034:13, :3049:13, :3064:13, :3079:13, :3094:13, :3109:13, :3124:13, :3139:13, :3154:13, :3169:13, :3184:13, :3199:13, :3214:13, :3229:13, :3244:13, :3259:13, :3274:13, :3289:13, :3304:13, :3319:13, :3334:13, :3349:13, :3364:13, :3379:13, :3394:13, :3409:13, :3424:13, :3439:13, :3454:13, :3469:13, :3484:13, :3499:13, :3514:13, :3529:13, :3544:13, :3559:13, :3574:13, :3589:13, :3604:13, :3619:13, :3634:13, :3649:13, :3664:13, :3679:13, :3694:13, :3709:13, :3724:13, :3739:13, :3754:13, :3769:13, :3784:13, :3799:13, :3814:13, :3829:13, :3844:13, :3847:13
  assign file_read_0_data = _T[file_read_0_addr];	// <stdin>:3846:13, :3849:5
  assign file_read_1_data = _T_0[file_read_1_addr];	// <stdin>:3848:13, :3849:5
endmodule

module code(	// <stdin>:3851:1
  input                                                        CLK, ASYNCRESET,
  input  [7:0]                                                 code_read_0_addr,
  input  struct packed {logic [31:0] data; logic [7:0] addr; } write_0,
  input                                                        write_0_en,
  output [31:0]                                                code_read_0_data);

  reg [31:0] Register_inst0;	// <stdin>:3859:10
  reg [31:0] Register_inst1;	// <stdin>:3875:11
  reg [31:0] Register_inst2;	// <stdin>:3890:11
  reg [31:0] Register_inst3;	// <stdin>:3905:11
  reg [31:0] Register_inst4;	// <stdin>:3920:11
  reg [31:0] Register_inst5;	// <stdin>:3935:11
  reg [31:0] Register_inst6;	// <stdin>:3950:11
  reg [31:0] Register_inst7;	// <stdin>:3965:11
  reg [31:0] Register_inst8;	// <stdin>:3980:11
  reg [31:0] Register_inst9;	// <stdin>:3995:11
  reg [31:0] Register_inst10;	// <stdin>:4010:11
  reg [31:0] Register_inst11;	// <stdin>:4025:11
  reg [31:0] Register_inst12;	// <stdin>:4040:11
  reg [31:0] Register_inst13;	// <stdin>:4055:12
  reg [31:0] Register_inst14;	// <stdin>:4070:12
  reg [31:0] Register_inst15;	// <stdin>:4085:12
  reg [31:0] Register_inst16;	// <stdin>:4100:12
  reg [31:0] Register_inst17;	// <stdin>:4115:12
  reg [31:0] Register_inst18;	// <stdin>:4130:12
  reg [31:0] Register_inst19;	// <stdin>:4145:12
  reg [31:0] Register_inst20;	// <stdin>:4160:12
  reg [31:0] Register_inst21;	// <stdin>:4175:12
  reg [31:0] Register_inst22;	// <stdin>:4190:12
  reg [31:0] Register_inst23;	// <stdin>:4205:12
  reg [31:0] Register_inst24;	// <stdin>:4220:12
  reg [31:0] Register_inst25;	// <stdin>:4235:12
  reg [31:0] Register_inst26;	// <stdin>:4250:12
  reg [31:0] Register_inst27;	// <stdin>:4265:12
  reg [31:0] Register_inst28;	// <stdin>:4280:12
  reg [31:0] Register_inst29;	// <stdin>:4295:12
  reg [31:0] Register_inst30;	// <stdin>:4310:12
  reg [31:0] Register_inst31;	// <stdin>:4325:12
  reg [31:0] Register_inst32;	// <stdin>:4340:12
  reg [31:0] Register_inst33;	// <stdin>:4355:12
  reg [31:0] Register_inst34;	// <stdin>:4370:12
  reg [31:0] Register_inst35;	// <stdin>:4385:12
  reg [31:0] Register_inst36;	// <stdin>:4400:12
  reg [31:0] Register_inst37;	// <stdin>:4415:12
  reg [31:0] Register_inst38;	// <stdin>:4430:12
  reg [31:0] Register_inst39;	// <stdin>:4445:12
  reg [31:0] Register_inst40;	// <stdin>:4460:12
  reg [31:0] Register_inst41;	// <stdin>:4475:12
  reg [31:0] Register_inst42;	// <stdin>:4490:12
  reg [31:0] Register_inst43;	// <stdin>:4505:12
  reg [31:0] Register_inst44;	// <stdin>:4520:12
  reg [31:0] Register_inst45;	// <stdin>:4535:12
  reg [31:0] Register_inst46;	// <stdin>:4550:12
  reg [31:0] Register_inst47;	// <stdin>:4565:12
  reg [31:0] Register_inst48;	// <stdin>:4580:12
  reg [31:0] Register_inst49;	// <stdin>:4595:12
  reg [31:0] Register_inst50;	// <stdin>:4610:12
  reg [31:0] Register_inst51;	// <stdin>:4625:12
  reg [31:0] Register_inst52;	// <stdin>:4640:12
  reg [31:0] Register_inst53;	// <stdin>:4655:12
  reg [31:0] Register_inst54;	// <stdin>:4670:12
  reg [31:0] Register_inst55;	// <stdin>:4685:12
  reg [31:0] Register_inst56;	// <stdin>:4700:12
  reg [31:0] Register_inst57;	// <stdin>:4715:12
  reg [31:0] Register_inst58;	// <stdin>:4730:12
  reg [31:0] Register_inst59;	// <stdin>:4745:12
  reg [31:0] Register_inst60;	// <stdin>:4760:12
  reg [31:0] Register_inst61;	// <stdin>:4775:12
  reg [31:0] Register_inst62;	// <stdin>:4790:12
  reg [31:0] Register_inst63;	// <stdin>:4805:12
  reg [31:0] Register_inst64;	// <stdin>:4820:12
  reg [31:0] Register_inst65;	// <stdin>:4835:12
  reg [31:0] Register_inst66;	// <stdin>:4850:12
  reg [31:0] Register_inst67;	// <stdin>:4865:12
  reg [31:0] Register_inst68;	// <stdin>:4880:12
  reg [31:0] Register_inst69;	// <stdin>:4895:12
  reg [31:0] Register_inst70;	// <stdin>:4910:12
  reg [31:0] Register_inst71;	// <stdin>:4925:12
  reg [31:0] Register_inst72;	// <stdin>:4940:12
  reg [31:0] Register_inst73;	// <stdin>:4955:12
  reg [31:0] Register_inst74;	// <stdin>:4970:12
  reg [31:0] Register_inst75;	// <stdin>:4985:12
  reg [31:0] Register_inst76;	// <stdin>:5000:12
  reg [31:0] Register_inst77;	// <stdin>:5015:12
  reg [31:0] Register_inst78;	// <stdin>:5030:12
  reg [31:0] Register_inst79;	// <stdin>:5045:12
  reg [31:0] Register_inst80;	// <stdin>:5060:12
  reg [31:0] Register_inst81;	// <stdin>:5075:12
  reg [31:0] Register_inst82;	// <stdin>:5090:12
  reg [31:0] Register_inst83;	// <stdin>:5105:12
  reg [31:0] Register_inst84;	// <stdin>:5120:12
  reg [31:0] Register_inst85;	// <stdin>:5135:12
  reg [31:0] Register_inst86;	// <stdin>:5150:12
  reg [31:0] Register_inst87;	// <stdin>:5165:12
  reg [31:0] Register_inst88;	// <stdin>:5180:12
  reg [31:0] Register_inst89;	// <stdin>:5195:12
  reg [31:0] Register_inst90;	// <stdin>:5210:12
  reg [31:0] Register_inst91;	// <stdin>:5225:12
  reg [31:0] Register_inst92;	// <stdin>:5240:12
  reg [31:0] Register_inst93;	// <stdin>:5255:12
  reg [31:0] Register_inst94;	// <stdin>:5270:12
  reg [31:0] Register_inst95;	// <stdin>:5285:12
  reg [31:0] Register_inst96;	// <stdin>:5300:12
  reg [31:0] Register_inst97;	// <stdin>:5315:12
  reg [31:0] Register_inst98;	// <stdin>:5330:12
  reg [31:0] Register_inst99;	// <stdin>:5345:12
  reg [31:0] Register_inst100;	// <stdin>:5360:12
  reg [31:0] Register_inst101;	// <stdin>:5375:12
  reg [31:0] Register_inst102;	// <stdin>:5390:12
  reg [31:0] Register_inst103;	// <stdin>:5405:12
  reg [31:0] Register_inst104;	// <stdin>:5420:12
  reg [31:0] Register_inst105;	// <stdin>:5435:12
  reg [31:0] Register_inst106;	// <stdin>:5450:12
  reg [31:0] Register_inst107;	// <stdin>:5465:12
  reg [31:0] Register_inst108;	// <stdin>:5480:12
  reg [31:0] Register_inst109;	// <stdin>:5495:12
  reg [31:0] Register_inst110;	// <stdin>:5510:12
  reg [31:0] Register_inst111;	// <stdin>:5525:12
  reg [31:0] Register_inst112;	// <stdin>:5540:12
  reg [31:0] Register_inst113;	// <stdin>:5555:12
  reg [31:0] Register_inst114;	// <stdin>:5570:12
  reg [31:0] Register_inst115;	// <stdin>:5585:12
  reg [31:0] Register_inst116;	// <stdin>:5600:12
  reg [31:0] Register_inst117;	// <stdin>:5615:12
  reg [31:0] Register_inst118;	// <stdin>:5630:12
  reg [31:0] Register_inst119;	// <stdin>:5645:12
  reg [31:0] Register_inst120;	// <stdin>:5660:12
  reg [31:0] Register_inst121;	// <stdin>:5675:12
  reg [31:0] Register_inst122;	// <stdin>:5690:12
  reg [31:0] Register_inst123;	// <stdin>:5705:12
  reg [31:0] Register_inst124;	// <stdin>:5720:12
  reg [31:0] Register_inst125;	// <stdin>:5735:12
  reg [31:0] Register_inst126;	// <stdin>:5750:12
  reg [31:0] Register_inst127;	// <stdin>:5765:12
  reg [31:0] Register_inst128;	// <stdin>:5780:12
  reg [31:0] Register_inst129;	// <stdin>:5795:12
  reg [31:0] Register_inst130;	// <stdin>:5810:12
  reg [31:0] Register_inst131;	// <stdin>:5825:12
  reg [31:0] Register_inst132;	// <stdin>:5840:12
  reg [31:0] Register_inst133;	// <stdin>:5855:12
  reg [31:0] Register_inst134;	// <stdin>:5870:12
  reg [31:0] Register_inst135;	// <stdin>:5885:12
  reg [31:0] Register_inst136;	// <stdin>:5900:12
  reg [31:0] Register_inst137;	// <stdin>:5915:12
  reg [31:0] Register_inst138;	// <stdin>:5930:12
  reg [31:0] Register_inst139;	// <stdin>:5945:12
  reg [31:0] Register_inst140;	// <stdin>:5960:12
  reg [31:0] Register_inst141;	// <stdin>:5975:12
  reg [31:0] Register_inst142;	// <stdin>:5990:13
  reg [31:0] Register_inst143;	// <stdin>:6005:13
  reg [31:0] Register_inst144;	// <stdin>:6020:13
  reg [31:0] Register_inst145;	// <stdin>:6035:13
  reg [31:0] Register_inst146;	// <stdin>:6050:13
  reg [31:0] Register_inst147;	// <stdin>:6065:13
  reg [31:0] Register_inst148;	// <stdin>:6080:13
  reg [31:0] Register_inst149;	// <stdin>:6095:13
  reg [31:0] Register_inst150;	// <stdin>:6110:13
  reg [31:0] Register_inst151;	// <stdin>:6125:13
  reg [31:0] Register_inst152;	// <stdin>:6140:13
  reg [31:0] Register_inst153;	// <stdin>:6155:13
  reg [31:0] Register_inst154;	// <stdin>:6170:13
  reg [31:0] Register_inst155;	// <stdin>:6185:13
  reg [31:0] Register_inst156;	// <stdin>:6200:13
  reg [31:0] Register_inst157;	// <stdin>:6215:13
  reg [31:0] Register_inst158;	// <stdin>:6230:13
  reg [31:0] Register_inst159;	// <stdin>:6245:13
  reg [31:0] Register_inst160;	// <stdin>:6260:13
  reg [31:0] Register_inst161;	// <stdin>:6275:13
  reg [31:0] Register_inst162;	// <stdin>:6290:13
  reg [31:0] Register_inst163;	// <stdin>:6305:13
  reg [31:0] Register_inst164;	// <stdin>:6320:13
  reg [31:0] Register_inst165;	// <stdin>:6335:13
  reg [31:0] Register_inst166;	// <stdin>:6350:13
  reg [31:0] Register_inst167;	// <stdin>:6365:13
  reg [31:0] Register_inst168;	// <stdin>:6380:13
  reg [31:0] Register_inst169;	// <stdin>:6395:13
  reg [31:0] Register_inst170;	// <stdin>:6410:13
  reg [31:0] Register_inst171;	// <stdin>:6425:13
  reg [31:0] Register_inst172;	// <stdin>:6440:13
  reg [31:0] Register_inst173;	// <stdin>:6455:13
  reg [31:0] Register_inst174;	// <stdin>:6470:13
  reg [31:0] Register_inst175;	// <stdin>:6485:13
  reg [31:0] Register_inst176;	// <stdin>:6500:13
  reg [31:0] Register_inst177;	// <stdin>:6515:13
  reg [31:0] Register_inst178;	// <stdin>:6530:13
  reg [31:0] Register_inst179;	// <stdin>:6545:13
  reg [31:0] Register_inst180;	// <stdin>:6560:13
  reg [31:0] Register_inst181;	// <stdin>:6575:13
  reg [31:0] Register_inst182;	// <stdin>:6590:13
  reg [31:0] Register_inst183;	// <stdin>:6605:13
  reg [31:0] Register_inst184;	// <stdin>:6620:13
  reg [31:0] Register_inst185;	// <stdin>:6635:13
  reg [31:0] Register_inst186;	// <stdin>:6650:13
  reg [31:0] Register_inst187;	// <stdin>:6665:13
  reg [31:0] Register_inst188;	// <stdin>:6680:13
  reg [31:0] Register_inst189;	// <stdin>:6695:13
  reg [31:0] Register_inst190;	// <stdin>:6710:13
  reg [31:0] Register_inst191;	// <stdin>:6725:13
  reg [31:0] Register_inst192;	// <stdin>:6740:13
  reg [31:0] Register_inst193;	// <stdin>:6755:13
  reg [31:0] Register_inst194;	// <stdin>:6770:13
  reg [31:0] Register_inst195;	// <stdin>:6785:13
  reg [31:0] Register_inst196;	// <stdin>:6800:13
  reg [31:0] Register_inst197;	// <stdin>:6815:13
  reg [31:0] Register_inst198;	// <stdin>:6830:13
  reg [31:0] Register_inst199;	// <stdin>:6845:13
  reg [31:0] Register_inst200;	// <stdin>:6860:13
  reg [31:0] Register_inst201;	// <stdin>:6875:13
  reg [31:0] Register_inst202;	// <stdin>:6890:13
  reg [31:0] Register_inst203;	// <stdin>:6905:13
  reg [31:0] Register_inst204;	// <stdin>:6920:13
  reg [31:0] Register_inst205;	// <stdin>:6935:13
  reg [31:0] Register_inst206;	// <stdin>:6950:13
  reg [31:0] Register_inst207;	// <stdin>:6965:13
  reg [31:0] Register_inst208;	// <stdin>:6980:13
  reg [31:0] Register_inst209;	// <stdin>:6995:13
  reg [31:0] Register_inst210;	// <stdin>:7010:13
  reg [31:0] Register_inst211;	// <stdin>:7025:13
  reg [31:0] Register_inst212;	// <stdin>:7040:13
  reg [31:0] Register_inst213;	// <stdin>:7055:13
  reg [31:0] Register_inst214;	// <stdin>:7070:13
  reg [31:0] Register_inst215;	// <stdin>:7085:13
  reg [31:0] Register_inst216;	// <stdin>:7100:13
  reg [31:0] Register_inst217;	// <stdin>:7115:13
  reg [31:0] Register_inst218;	// <stdin>:7130:13
  reg [31:0] Register_inst219;	// <stdin>:7145:13
  reg [31:0] Register_inst220;	// <stdin>:7160:13
  reg [31:0] Register_inst221;	// <stdin>:7175:13
  reg [31:0] Register_inst222;	// <stdin>:7190:13
  reg [31:0] Register_inst223;	// <stdin>:7205:13
  reg [31:0] Register_inst224;	// <stdin>:7220:13
  reg [31:0] Register_inst225;	// <stdin>:7235:13
  reg [31:0] Register_inst226;	// <stdin>:7250:13
  reg [31:0] Register_inst227;	// <stdin>:7265:13
  reg [31:0] Register_inst228;	// <stdin>:7280:13
  reg [31:0] Register_inst229;	// <stdin>:7295:13
  reg [31:0] Register_inst230;	// <stdin>:7310:13
  reg [31:0] Register_inst231;	// <stdin>:7325:13
  reg [31:0] Register_inst232;	// <stdin>:7340:13
  reg [31:0] Register_inst233;	// <stdin>:7355:13
  reg [31:0] Register_inst234;	// <stdin>:7370:13
  reg [31:0] Register_inst235;	// <stdin>:7385:13
  reg [31:0] Register_inst236;	// <stdin>:7400:13
  reg [31:0] Register_inst237;	// <stdin>:7415:13
  reg [31:0] Register_inst238;	// <stdin>:7430:13
  reg [31:0] Register_inst239;	// <stdin>:7445:13
  reg [31:0] Register_inst240;	// <stdin>:7460:13
  reg [31:0] Register_inst241;	// <stdin>:7475:13
  reg [31:0] Register_inst242;	// <stdin>:7490:13
  reg [31:0] Register_inst243;	// <stdin>:7505:13
  reg [31:0] Register_inst244;	// <stdin>:7520:13
  reg [31:0] Register_inst245;	// <stdin>:7535:13
  reg [31:0] Register_inst246;	// <stdin>:7550:13
  reg [31:0] Register_inst247;	// <stdin>:7565:13
  reg [31:0] Register_inst248;	// <stdin>:7580:13
  reg [31:0] Register_inst249;	// <stdin>:7595:13
  reg [31:0] Register_inst250;	// <stdin>:7610:13
  reg [31:0] Register_inst251;	// <stdin>:7625:13
  reg [31:0] Register_inst252;	// <stdin>:7640:13
  reg [31:0] Register_inst253;	// <stdin>:7655:13
  reg [31:0] Register_inst254;	// <stdin>:7670:13
  reg [31:0] Register_inst255;	// <stdin>:7685:13

  always_ff @(posedge CLK or posedge ASYNCRESET) begin	// <stdin>:7686:5
    if (ASYNCRESET) begin	// <stdin>:7686:5
      Register_inst0 <= 32'h0;	// <stdin>:3863:9, :3865:10
      Register_inst1 <= 32'h0;	// <stdin>:3865:10, :3879:9
      Register_inst2 <= 32'h0;	// <stdin>:3865:10, :3894:9
      Register_inst3 <= 32'h0;	// <stdin>:3865:10, :3909:9
      Register_inst4 <= 32'h0;	// <stdin>:3865:10, :3924:9
      Register_inst5 <= 32'h0;	// <stdin>:3865:10, :3939:9
      Register_inst6 <= 32'h0;	// <stdin>:3865:10, :3954:9
      Register_inst7 <= 32'h0;	// <stdin>:3865:10, :3969:9
      Register_inst8 <= 32'h0;	// <stdin>:3865:10, :3984:9
      Register_inst9 <= 32'h0;	// <stdin>:3865:10, :3999:9
      Register_inst10 <= 32'h0;	// <stdin>:3865:10, :4014:9
      Register_inst11 <= 32'h0;	// <stdin>:3865:10, :4029:9
      Register_inst12 <= 32'h0;	// <stdin>:3865:10, :4044:9
      Register_inst13 <= 32'h0;	// <stdin>:3865:10, :4059:9
      Register_inst14 <= 32'h0;	// <stdin>:3865:10, :4074:9
      Register_inst15 <= 32'h0;	// <stdin>:3865:10, :4089:9
      Register_inst16 <= 32'h0;	// <stdin>:3865:10, :4104:9
      Register_inst17 <= 32'h0;	// <stdin>:3865:10, :4119:9
      Register_inst18 <= 32'h0;	// <stdin>:3865:10, :4134:9
      Register_inst19 <= 32'h0;	// <stdin>:3865:10, :4149:9
      Register_inst20 <= 32'h0;	// <stdin>:3865:10, :4164:9
      Register_inst21 <= 32'h0;	// <stdin>:3865:10, :4179:9
      Register_inst22 <= 32'h0;	// <stdin>:3865:10, :4194:9
      Register_inst23 <= 32'h0;	// <stdin>:3865:10, :4209:9
      Register_inst24 <= 32'h0;	// <stdin>:3865:10, :4224:9
      Register_inst25 <= 32'h0;	// <stdin>:3865:10, :4239:9
      Register_inst26 <= 32'h0;	// <stdin>:3865:10, :4254:9
      Register_inst27 <= 32'h0;	// <stdin>:3865:10, :4269:9
      Register_inst28 <= 32'h0;	// <stdin>:3865:10, :4284:9
      Register_inst29 <= 32'h0;	// <stdin>:3865:10, :4299:9
      Register_inst30 <= 32'h0;	// <stdin>:3865:10, :4314:9
      Register_inst31 <= 32'h0;	// <stdin>:3865:10, :4329:9
      Register_inst32 <= 32'h0;	// <stdin>:3865:10, :4344:9
      Register_inst33 <= 32'h0;	// <stdin>:3865:10, :4359:9
      Register_inst34 <= 32'h0;	// <stdin>:3865:10, :4374:9
      Register_inst35 <= 32'h0;	// <stdin>:3865:10, :4389:9
      Register_inst36 <= 32'h0;	// <stdin>:3865:10, :4404:9
      Register_inst37 <= 32'h0;	// <stdin>:3865:10, :4419:9
      Register_inst38 <= 32'h0;	// <stdin>:3865:10, :4434:9
      Register_inst39 <= 32'h0;	// <stdin>:3865:10, :4449:9
      Register_inst40 <= 32'h0;	// <stdin>:3865:10, :4464:9
      Register_inst41 <= 32'h0;	// <stdin>:3865:10, :4479:9
      Register_inst42 <= 32'h0;	// <stdin>:3865:10, :4494:9
      Register_inst43 <= 32'h0;	// <stdin>:3865:10, :4509:9
      Register_inst44 <= 32'h0;	// <stdin>:3865:10, :4524:9
      Register_inst45 <= 32'h0;	// <stdin>:3865:10, :4539:9
      Register_inst46 <= 32'h0;	// <stdin>:3865:10, :4554:9
      Register_inst47 <= 32'h0;	// <stdin>:3865:10, :4569:9
      Register_inst48 <= 32'h0;	// <stdin>:3865:10, :4584:9
      Register_inst49 <= 32'h0;	// <stdin>:3865:10, :4599:9
      Register_inst50 <= 32'h0;	// <stdin>:3865:10, :4614:9
      Register_inst51 <= 32'h0;	// <stdin>:3865:10, :4629:9
      Register_inst52 <= 32'h0;	// <stdin>:3865:10, :4644:9
      Register_inst53 <= 32'h0;	// <stdin>:3865:10, :4659:9
      Register_inst54 <= 32'h0;	// <stdin>:3865:10, :4674:9
      Register_inst55 <= 32'h0;	// <stdin>:3865:10, :4689:9
      Register_inst56 <= 32'h0;	// <stdin>:3865:10, :4704:9
      Register_inst57 <= 32'h0;	// <stdin>:3865:10, :4719:9
      Register_inst58 <= 32'h0;	// <stdin>:3865:10, :4734:9
      Register_inst59 <= 32'h0;	// <stdin>:3865:10, :4749:9
      Register_inst60 <= 32'h0;	// <stdin>:3865:10, :4764:9
      Register_inst61 <= 32'h0;	// <stdin>:3865:10, :4779:9
      Register_inst62 <= 32'h0;	// <stdin>:3865:10, :4794:9
      Register_inst63 <= 32'h0;	// <stdin>:3865:10, :4809:9
      Register_inst64 <= 32'h0;	// <stdin>:3865:10, :4824:9
      Register_inst65 <= 32'h0;	// <stdin>:3865:10, :4839:9
      Register_inst66 <= 32'h0;	// <stdin>:3865:10, :4854:9
      Register_inst67 <= 32'h0;	// <stdin>:3865:10, :4869:9
      Register_inst68 <= 32'h0;	// <stdin>:3865:10, :4884:9
      Register_inst69 <= 32'h0;	// <stdin>:3865:10, :4899:9
      Register_inst70 <= 32'h0;	// <stdin>:3865:10, :4914:9
      Register_inst71 <= 32'h0;	// <stdin>:3865:10, :4929:9
      Register_inst72 <= 32'h0;	// <stdin>:3865:10, :4944:9
      Register_inst73 <= 32'h0;	// <stdin>:3865:10, :4959:9
      Register_inst74 <= 32'h0;	// <stdin>:3865:10, :4974:9
      Register_inst75 <= 32'h0;	// <stdin>:3865:10, :4989:9
      Register_inst76 <= 32'h0;	// <stdin>:3865:10, :5004:9
      Register_inst77 <= 32'h0;	// <stdin>:3865:10, :5019:9
      Register_inst78 <= 32'h0;	// <stdin>:3865:10, :5034:9
      Register_inst79 <= 32'h0;	// <stdin>:3865:10, :5049:9
      Register_inst80 <= 32'h0;	// <stdin>:3865:10, :5064:9
      Register_inst81 <= 32'h0;	// <stdin>:3865:10, :5079:9
      Register_inst82 <= 32'h0;	// <stdin>:3865:10, :5094:9
      Register_inst83 <= 32'h0;	// <stdin>:3865:10, :5109:9
      Register_inst84 <= 32'h0;	// <stdin>:3865:10, :5124:9
      Register_inst85 <= 32'h0;	// <stdin>:3865:10, :5139:9
      Register_inst86 <= 32'h0;	// <stdin>:3865:10, :5154:9
      Register_inst87 <= 32'h0;	// <stdin>:3865:10, :5169:9
      Register_inst88 <= 32'h0;	// <stdin>:3865:10, :5184:9
      Register_inst89 <= 32'h0;	// <stdin>:3865:10, :5199:9
      Register_inst90 <= 32'h0;	// <stdin>:3865:10, :5214:9
      Register_inst91 <= 32'h0;	// <stdin>:3865:10, :5229:9
      Register_inst92 <= 32'h0;	// <stdin>:3865:10, :5244:9
      Register_inst93 <= 32'h0;	// <stdin>:3865:10, :5259:9
      Register_inst94 <= 32'h0;	// <stdin>:3865:10, :5274:9
      Register_inst95 <= 32'h0;	// <stdin>:3865:10, :5289:9
      Register_inst96 <= 32'h0;	// <stdin>:3865:10, :5304:9
      Register_inst97 <= 32'h0;	// <stdin>:3865:10, :5319:9
      Register_inst98 <= 32'h0;	// <stdin>:3865:10, :5334:9
      Register_inst99 <= 32'h0;	// <stdin>:3865:10, :5349:9
      Register_inst100 <= 32'h0;	// <stdin>:3865:10, :5364:9
      Register_inst101 <= 32'h0;	// <stdin>:3865:10, :5379:9
      Register_inst102 <= 32'h0;	// <stdin>:3865:10, :5394:9
      Register_inst103 <= 32'h0;	// <stdin>:3865:10, :5409:9
      Register_inst104 <= 32'h0;	// <stdin>:3865:10, :5424:9
      Register_inst105 <= 32'h0;	// <stdin>:3865:10, :5439:9
      Register_inst106 <= 32'h0;	// <stdin>:3865:10, :5454:9
      Register_inst107 <= 32'h0;	// <stdin>:3865:10, :5469:9
      Register_inst108 <= 32'h0;	// <stdin>:3865:10, :5484:9
      Register_inst109 <= 32'h0;	// <stdin>:3865:10, :5499:9
      Register_inst110 <= 32'h0;	// <stdin>:3865:10, :5514:9
      Register_inst111 <= 32'h0;	// <stdin>:3865:10, :5529:9
      Register_inst112 <= 32'h0;	// <stdin>:3865:10, :5544:9
      Register_inst113 <= 32'h0;	// <stdin>:3865:10, :5559:9
      Register_inst114 <= 32'h0;	// <stdin>:3865:10, :5574:9
      Register_inst115 <= 32'h0;	// <stdin>:3865:10, :5589:9
      Register_inst116 <= 32'h0;	// <stdin>:3865:10, :5604:9
      Register_inst117 <= 32'h0;	// <stdin>:3865:10, :5619:9
      Register_inst118 <= 32'h0;	// <stdin>:3865:10, :5634:9
      Register_inst119 <= 32'h0;	// <stdin>:3865:10, :5649:9
      Register_inst120 <= 32'h0;	// <stdin>:3865:10, :5664:9
      Register_inst121 <= 32'h0;	// <stdin>:3865:10, :5679:9
      Register_inst122 <= 32'h0;	// <stdin>:3865:10, :5694:9
      Register_inst123 <= 32'h0;	// <stdin>:3865:10, :5709:9
      Register_inst124 <= 32'h0;	// <stdin>:3865:10, :5724:9
      Register_inst125 <= 32'h0;	// <stdin>:3865:10, :5739:9
      Register_inst126 <= 32'h0;	// <stdin>:3865:10, :5754:9
      Register_inst127 <= 32'h0;	// <stdin>:3865:10, :5769:9
      Register_inst128 <= 32'h0;	// <stdin>:3865:10, :5784:9
      Register_inst129 <= 32'h0;	// <stdin>:3865:10, :5799:9
      Register_inst130 <= 32'h0;	// <stdin>:3865:10, :5814:9
      Register_inst131 <= 32'h0;	// <stdin>:3865:10, :5829:9
      Register_inst132 <= 32'h0;	// <stdin>:3865:10, :5844:9
      Register_inst133 <= 32'h0;	// <stdin>:3865:10, :5859:9
      Register_inst134 <= 32'h0;	// <stdin>:3865:10, :5874:9
      Register_inst135 <= 32'h0;	// <stdin>:3865:10, :5889:9
      Register_inst136 <= 32'h0;	// <stdin>:3865:10, :5904:9
      Register_inst137 <= 32'h0;	// <stdin>:3865:10, :5919:9
      Register_inst138 <= 32'h0;	// <stdin>:3865:10, :5934:9
      Register_inst139 <= 32'h0;	// <stdin>:3865:10, :5949:9
      Register_inst140 <= 32'h0;	// <stdin>:3865:10, :5964:9
      Register_inst141 <= 32'h0;	// <stdin>:3865:10, :5979:9
      Register_inst142 <= 32'h0;	// <stdin>:3865:10, :5994:9
      Register_inst143 <= 32'h0;	// <stdin>:3865:10, :6009:9
      Register_inst144 <= 32'h0;	// <stdin>:3865:10, :6024:9
      Register_inst145 <= 32'h0;	// <stdin>:3865:10, :6039:9
      Register_inst146 <= 32'h0;	// <stdin>:3865:10, :6054:9
      Register_inst147 <= 32'h0;	// <stdin>:3865:10, :6069:9
      Register_inst148 <= 32'h0;	// <stdin>:3865:10, :6084:9
      Register_inst149 <= 32'h0;	// <stdin>:3865:10, :6099:9
      Register_inst150 <= 32'h0;	// <stdin>:3865:10, :6114:9
      Register_inst151 <= 32'h0;	// <stdin>:3865:10, :6129:9
      Register_inst152 <= 32'h0;	// <stdin>:3865:10, :6144:9
      Register_inst153 <= 32'h0;	// <stdin>:3865:10, :6159:9
      Register_inst154 <= 32'h0;	// <stdin>:3865:10, :6174:9
      Register_inst155 <= 32'h0;	// <stdin>:3865:10, :6189:9
      Register_inst156 <= 32'h0;	// <stdin>:3865:10, :6204:9
      Register_inst157 <= 32'h0;	// <stdin>:3865:10, :6219:9
      Register_inst158 <= 32'h0;	// <stdin>:3865:10, :6234:9
      Register_inst159 <= 32'h0;	// <stdin>:3865:10, :6249:9
      Register_inst160 <= 32'h0;	// <stdin>:3865:10, :6264:9
      Register_inst161 <= 32'h0;	// <stdin>:3865:10, :6279:9
      Register_inst162 <= 32'h0;	// <stdin>:3865:10, :6294:9
      Register_inst163 <= 32'h0;	// <stdin>:3865:10, :6309:9
      Register_inst164 <= 32'h0;	// <stdin>:3865:10, :6324:9
      Register_inst165 <= 32'h0;	// <stdin>:3865:10, :6339:9
      Register_inst166 <= 32'h0;	// <stdin>:3865:10, :6354:9
      Register_inst167 <= 32'h0;	// <stdin>:3865:10, :6369:9
      Register_inst168 <= 32'h0;	// <stdin>:3865:10, :6384:9
      Register_inst169 <= 32'h0;	// <stdin>:3865:10, :6399:9
      Register_inst170 <= 32'h0;	// <stdin>:3865:10, :6414:9
      Register_inst171 <= 32'h0;	// <stdin>:3865:10, :6429:9
      Register_inst172 <= 32'h0;	// <stdin>:3865:10, :6444:9
      Register_inst173 <= 32'h0;	// <stdin>:3865:10, :6459:9
      Register_inst174 <= 32'h0;	// <stdin>:3865:10, :6474:9
      Register_inst175 <= 32'h0;	// <stdin>:3865:10, :6489:9
      Register_inst176 <= 32'h0;	// <stdin>:3865:10, :6504:9
      Register_inst177 <= 32'h0;	// <stdin>:3865:10, :6519:9
      Register_inst178 <= 32'h0;	// <stdin>:3865:10, :6534:9
      Register_inst179 <= 32'h0;	// <stdin>:3865:10, :6549:9
      Register_inst180 <= 32'h0;	// <stdin>:3865:10, :6564:9
      Register_inst181 <= 32'h0;	// <stdin>:3865:10, :6579:9
      Register_inst182 <= 32'h0;	// <stdin>:3865:10, :6594:9
      Register_inst183 <= 32'h0;	// <stdin>:3865:10, :6609:9
      Register_inst184 <= 32'h0;	// <stdin>:3865:10, :6624:9
      Register_inst185 <= 32'h0;	// <stdin>:3865:10, :6639:9
      Register_inst186 <= 32'h0;	// <stdin>:3865:10, :6654:9
      Register_inst187 <= 32'h0;	// <stdin>:3865:10, :6669:9
      Register_inst188 <= 32'h0;	// <stdin>:3865:10, :6684:9
      Register_inst189 <= 32'h0;	// <stdin>:3865:10, :6699:9
      Register_inst190 <= 32'h0;	// <stdin>:3865:10, :6714:9
      Register_inst191 <= 32'h0;	// <stdin>:3865:10, :6729:9
      Register_inst192 <= 32'h0;	// <stdin>:3865:10, :6744:9
      Register_inst193 <= 32'h0;	// <stdin>:3865:10, :6759:9
      Register_inst194 <= 32'h0;	// <stdin>:3865:10, :6774:9
      Register_inst195 <= 32'h0;	// <stdin>:3865:10, :6789:9
      Register_inst196 <= 32'h0;	// <stdin>:3865:10, :6804:9
      Register_inst197 <= 32'h0;	// <stdin>:3865:10, :6819:9
      Register_inst198 <= 32'h0;	// <stdin>:3865:10, :6834:9
      Register_inst199 <= 32'h0;	// <stdin>:3865:10, :6849:9
      Register_inst200 <= 32'h0;	// <stdin>:3865:10, :6864:9
      Register_inst201 <= 32'h0;	// <stdin>:3865:10, :6879:9
      Register_inst202 <= 32'h0;	// <stdin>:3865:10, :6894:9
      Register_inst203 <= 32'h0;	// <stdin>:3865:10, :6909:9
      Register_inst204 <= 32'h0;	// <stdin>:3865:10, :6924:9
      Register_inst205 <= 32'h0;	// <stdin>:3865:10, :6939:9
      Register_inst206 <= 32'h0;	// <stdin>:3865:10, :6954:9
      Register_inst207 <= 32'h0;	// <stdin>:3865:10, :6969:9
      Register_inst208 <= 32'h0;	// <stdin>:3865:10, :6984:9
      Register_inst209 <= 32'h0;	// <stdin>:3865:10, :6999:9
      Register_inst210 <= 32'h0;	// <stdin>:3865:10, :7014:9
      Register_inst211 <= 32'h0;	// <stdin>:3865:10, :7029:9
      Register_inst212 <= 32'h0;	// <stdin>:3865:10, :7044:9
      Register_inst213 <= 32'h0;	// <stdin>:3865:10, :7059:9
      Register_inst214 <= 32'h0;	// <stdin>:3865:10, :7074:9
      Register_inst215 <= 32'h0;	// <stdin>:3865:10, :7089:9
      Register_inst216 <= 32'h0;	// <stdin>:3865:10, :7104:9
      Register_inst217 <= 32'h0;	// <stdin>:3865:10, :7119:9
      Register_inst218 <= 32'h0;	// <stdin>:3865:10, :7134:9
      Register_inst219 <= 32'h0;	// <stdin>:3865:10, :7149:9
      Register_inst220 <= 32'h0;	// <stdin>:3865:10, :7164:9
      Register_inst221 <= 32'h0;	// <stdin>:3865:10, :7179:9
      Register_inst222 <= 32'h0;	// <stdin>:3865:10, :7194:9
      Register_inst223 <= 32'h0;	// <stdin>:3865:10, :7209:9
      Register_inst224 <= 32'h0;	// <stdin>:3865:10, :7224:9
      Register_inst225 <= 32'h0;	// <stdin>:3865:10, :7239:9
      Register_inst226 <= 32'h0;	// <stdin>:3865:10, :7254:9
      Register_inst227 <= 32'h0;	// <stdin>:3865:10, :7269:9
      Register_inst228 <= 32'h0;	// <stdin>:3865:10, :7284:9
      Register_inst229 <= 32'h0;	// <stdin>:3865:10, :7299:9
      Register_inst230 <= 32'h0;	// <stdin>:3865:10, :7314:9
      Register_inst231 <= 32'h0;	// <stdin>:3865:10, :7329:9
      Register_inst232 <= 32'h0;	// <stdin>:3865:10, :7344:9
      Register_inst233 <= 32'h0;	// <stdin>:3865:10, :7359:9
      Register_inst234 <= 32'h0;	// <stdin>:3865:10, :7374:9
      Register_inst235 <= 32'h0;	// <stdin>:3865:10, :7389:9
      Register_inst236 <= 32'h0;	// <stdin>:3865:10, :7404:9
      Register_inst237 <= 32'h0;	// <stdin>:3865:10, :7419:9
      Register_inst238 <= 32'h0;	// <stdin>:3865:10, :7434:9
      Register_inst239 <= 32'h0;	// <stdin>:3865:10, :7449:9
      Register_inst240 <= 32'h0;	// <stdin>:3865:10, :7464:9
      Register_inst241 <= 32'h0;	// <stdin>:3865:10, :7479:9
      Register_inst242 <= 32'h0;	// <stdin>:3865:10, :7494:9
      Register_inst243 <= 32'h0;	// <stdin>:3865:10, :7509:9
      Register_inst244 <= 32'h0;	// <stdin>:3865:10, :7524:9
      Register_inst245 <= 32'h0;	// <stdin>:3865:10, :7539:9
      Register_inst246 <= 32'h0;	// <stdin>:3865:10, :7554:9
      Register_inst247 <= 32'h0;	// <stdin>:3865:10, :7569:9
      Register_inst248 <= 32'h0;	// <stdin>:3865:10, :7584:9
      Register_inst249 <= 32'h0;	// <stdin>:3865:10, :7599:9
      Register_inst250 <= 32'h0;	// <stdin>:3865:10, :7614:9
      Register_inst251 <= 32'h0;	// <stdin>:3865:10, :7629:9
      Register_inst252 <= 32'h0;	// <stdin>:3865:10, :7644:9
      Register_inst253 <= 32'h0;	// <stdin>:3865:10, :7659:9
      Register_inst254 <= 32'h0;	// <stdin>:3865:10, :7674:9
      Register_inst255 <= 32'h0;	// <stdin>:3865:10, :7689:9
    end
    else begin	// <stdin>:7686:5
      automatic logic [31:0]      _T_0 = write_0.data;	// <stdin>:3852:10
      automatic logic [7:0]       _T_1 = write_0.addr;	// <stdin>:3853:10
      automatic logic [1:0][31:0] _T_2 = {{Register_inst0}, {_T_0}};	// <stdin>:3857:10, :3869:10
      automatic logic [1:0][31:0] _T_3 = {{Register_inst1}, {_T_0}};	// <stdin>:3873:11, :3884:11
      automatic logic [1:0][31:0] _T_4 = {{Register_inst2}, {_T_0}};	// <stdin>:3888:11, :3899:11
      automatic logic [1:0][31:0] _T_5 = {{Register_inst3}, {_T_0}};	// <stdin>:3903:11, :3914:11
      automatic logic [1:0][31:0] _T_6 = {{Register_inst4}, {_T_0}};	// <stdin>:3918:11, :3929:11
      automatic logic [1:0][31:0] _T_7 = {{Register_inst5}, {_T_0}};	// <stdin>:3933:11, :3944:11
      automatic logic [1:0][31:0] _T_8 = {{Register_inst6}, {_T_0}};	// <stdin>:3948:11, :3959:11
      automatic logic [1:0][31:0] _T_9 = {{Register_inst7}, {_T_0}};	// <stdin>:3963:11, :3974:11
      automatic logic [1:0][31:0] _T_10 = {{Register_inst8}, {_T_0}};	// <stdin>:3978:11, :3989:11
      automatic logic [1:0][31:0] _T_11 = {{Register_inst9}, {_T_0}};	// <stdin>:3993:11, :4004:11
      automatic logic [1:0][31:0] _T_12 = {{Register_inst10}, {_T_0}};	// <stdin>:4008:11, :4019:11
      automatic logic [1:0][31:0] _T_13 = {{Register_inst11}, {_T_0}};	// <stdin>:4023:11, :4034:11
      automatic logic [1:0][31:0] _T_14 = {{Register_inst12}, {_T_0}};	// <stdin>:4038:11, :4049:11
      automatic logic [1:0][31:0] _T_15 = {{Register_inst13}, {_T_0}};	// <stdin>:4053:11, :4064:11
      automatic logic [1:0][31:0] _T_16 = {{Register_inst14}, {_T_0}};	// <stdin>:4068:12, :4079:12
      automatic logic [1:0][31:0] _T_17 = {{Register_inst15}, {_T_0}};	// <stdin>:4083:12, :4094:12
      automatic logic [1:0][31:0] _T_18 = {{Register_inst16}, {_T_0}};	// <stdin>:4098:12, :4109:12
      automatic logic [1:0][31:0] _T_19 = {{Register_inst17}, {_T_0}};	// <stdin>:4113:12, :4124:12
      automatic logic [1:0][31:0] _T_20 = {{Register_inst18}, {_T_0}};	// <stdin>:4128:12, :4139:12
      automatic logic [1:0][31:0] _T_21 = {{Register_inst19}, {_T_0}};	// <stdin>:4143:12, :4154:12
      automatic logic [1:0][31:0] _T_22 = {{Register_inst20}, {_T_0}};	// <stdin>:4158:12, :4169:12
      automatic logic [1:0][31:0] _T_23 = {{Register_inst21}, {_T_0}};	// <stdin>:4173:12, :4184:12
      automatic logic [1:0][31:0] _T_24 = {{Register_inst22}, {_T_0}};	// <stdin>:4188:12, :4199:12
      automatic logic [1:0][31:0] _T_25 = {{Register_inst23}, {_T_0}};	// <stdin>:4203:12, :4214:12
      automatic logic [1:0][31:0] _T_26 = {{Register_inst24}, {_T_0}};	// <stdin>:4218:12, :4229:12
      automatic logic [1:0][31:0] _T_27 = {{Register_inst25}, {_T_0}};	// <stdin>:4233:12, :4244:12
      automatic logic [1:0][31:0] _T_28 = {{Register_inst26}, {_T_0}};	// <stdin>:4248:12, :4259:12
      automatic logic [1:0][31:0] _T_29 = {{Register_inst27}, {_T_0}};	// <stdin>:4263:12, :4274:12
      automatic logic [1:0][31:0] _T_30 = {{Register_inst28}, {_T_0}};	// <stdin>:4278:12, :4289:12
      automatic logic [1:0][31:0] _T_31 = {{Register_inst29}, {_T_0}};	// <stdin>:4293:12, :4304:12
      automatic logic [1:0][31:0] _T_32 = {{Register_inst30}, {_T_0}};	// <stdin>:4308:12, :4319:12
      automatic logic [1:0][31:0] _T_33 = {{Register_inst31}, {_T_0}};	// <stdin>:4323:12, :4334:12
      automatic logic [1:0][31:0] _T_34 = {{Register_inst32}, {_T_0}};	// <stdin>:4338:12, :4349:12
      automatic logic [1:0][31:0] _T_35 = {{Register_inst33}, {_T_0}};	// <stdin>:4353:12, :4364:12
      automatic logic [1:0][31:0] _T_36 = {{Register_inst34}, {_T_0}};	// <stdin>:4368:12, :4379:12
      automatic logic [1:0][31:0] _T_37 = {{Register_inst35}, {_T_0}};	// <stdin>:4383:12, :4394:12
      automatic logic [1:0][31:0] _T_38 = {{Register_inst36}, {_T_0}};	// <stdin>:4398:12, :4409:12
      automatic logic [1:0][31:0] _T_39 = {{Register_inst37}, {_T_0}};	// <stdin>:4413:12, :4424:12
      automatic logic [1:0][31:0] _T_40 = {{Register_inst38}, {_T_0}};	// <stdin>:4428:12, :4439:12
      automatic logic [1:0][31:0] _T_41 = {{Register_inst39}, {_T_0}};	// <stdin>:4443:12, :4454:12
      automatic logic [1:0][31:0] _T_42 = {{Register_inst40}, {_T_0}};	// <stdin>:4458:12, :4469:12
      automatic logic [1:0][31:0] _T_43 = {{Register_inst41}, {_T_0}};	// <stdin>:4473:12, :4484:12
      automatic logic [1:0][31:0] _T_44 = {{Register_inst42}, {_T_0}};	// <stdin>:4488:12, :4499:12
      automatic logic [1:0][31:0] _T_45 = {{Register_inst43}, {_T_0}};	// <stdin>:4503:12, :4514:12
      automatic logic [1:0][31:0] _T_46 = {{Register_inst44}, {_T_0}};	// <stdin>:4518:12, :4529:12
      automatic logic [1:0][31:0] _T_47 = {{Register_inst45}, {_T_0}};	// <stdin>:4533:12, :4544:12
      automatic logic [1:0][31:0] _T_48 = {{Register_inst46}, {_T_0}};	// <stdin>:4548:12, :4559:12
      automatic logic [1:0][31:0] _T_49 = {{Register_inst47}, {_T_0}};	// <stdin>:4563:12, :4574:12
      automatic logic [1:0][31:0] _T_50 = {{Register_inst48}, {_T_0}};	// <stdin>:4578:12, :4589:12
      automatic logic [1:0][31:0] _T_51 = {{Register_inst49}, {_T_0}};	// <stdin>:4593:12, :4604:12
      automatic logic [1:0][31:0] _T_52 = {{Register_inst50}, {_T_0}};	// <stdin>:4608:12, :4619:12
      automatic logic [1:0][31:0] _T_53 = {{Register_inst51}, {_T_0}};	// <stdin>:4623:12, :4634:12
      automatic logic [1:0][31:0] _T_54 = {{Register_inst52}, {_T_0}};	// <stdin>:4638:12, :4649:12
      automatic logic [1:0][31:0] _T_55 = {{Register_inst53}, {_T_0}};	// <stdin>:4653:12, :4664:12
      automatic logic [1:0][31:0] _T_56 = {{Register_inst54}, {_T_0}};	// <stdin>:4668:12, :4679:12
      automatic logic [1:0][31:0] _T_57 = {{Register_inst55}, {_T_0}};	// <stdin>:4683:12, :4694:12
      automatic logic [1:0][31:0] _T_58 = {{Register_inst56}, {_T_0}};	// <stdin>:4698:12, :4709:12
      automatic logic [1:0][31:0] _T_59 = {{Register_inst57}, {_T_0}};	// <stdin>:4713:12, :4724:12
      automatic logic [1:0][31:0] _T_60 = {{Register_inst58}, {_T_0}};	// <stdin>:4728:12, :4739:12
      automatic logic [1:0][31:0] _T_61 = {{Register_inst59}, {_T_0}};	// <stdin>:4743:12, :4754:12
      automatic logic [1:0][31:0] _T_62 = {{Register_inst60}, {_T_0}};	// <stdin>:4758:12, :4769:12
      automatic logic [1:0][31:0] _T_63 = {{Register_inst61}, {_T_0}};	// <stdin>:4773:12, :4784:12
      automatic logic [1:0][31:0] _T_64 = {{Register_inst62}, {_T_0}};	// <stdin>:4788:12, :4799:12
      automatic logic [1:0][31:0] _T_65 = {{Register_inst63}, {_T_0}};	// <stdin>:4803:12, :4814:12
      automatic logic [1:0][31:0] _T_66 = {{Register_inst64}, {_T_0}};	// <stdin>:4818:12, :4829:12
      automatic logic [1:0][31:0] _T_67 = {{Register_inst65}, {_T_0}};	// <stdin>:4833:12, :4844:12
      automatic logic [1:0][31:0] _T_68 = {{Register_inst66}, {_T_0}};	// <stdin>:4848:12, :4859:12
      automatic logic [1:0][31:0] _T_69 = {{Register_inst67}, {_T_0}};	// <stdin>:4863:12, :4874:12
      automatic logic [1:0][31:0] _T_70 = {{Register_inst68}, {_T_0}};	// <stdin>:4878:12, :4889:12
      automatic logic [1:0][31:0] _T_71 = {{Register_inst69}, {_T_0}};	// <stdin>:4893:12, :4904:12
      automatic logic [1:0][31:0] _T_72 = {{Register_inst70}, {_T_0}};	// <stdin>:4908:12, :4919:12
      automatic logic [1:0][31:0] _T_73 = {{Register_inst71}, {_T_0}};	// <stdin>:4923:12, :4934:12
      automatic logic [1:0][31:0] _T_74 = {{Register_inst72}, {_T_0}};	// <stdin>:4938:12, :4949:12
      automatic logic [1:0][31:0] _T_75 = {{Register_inst73}, {_T_0}};	// <stdin>:4953:12, :4964:12
      automatic logic [1:0][31:0] _T_76 = {{Register_inst74}, {_T_0}};	// <stdin>:4968:12, :4979:12
      automatic logic [1:0][31:0] _T_77 = {{Register_inst75}, {_T_0}};	// <stdin>:4983:12, :4994:12
      automatic logic [1:0][31:0] _T_78 = {{Register_inst76}, {_T_0}};	// <stdin>:4998:12, :5009:12
      automatic logic [1:0][31:0] _T_79 = {{Register_inst77}, {_T_0}};	// <stdin>:5013:12, :5024:12
      automatic logic [1:0][31:0] _T_80 = {{Register_inst78}, {_T_0}};	// <stdin>:5028:12, :5039:12
      automatic logic [1:0][31:0] _T_81 = {{Register_inst79}, {_T_0}};	// <stdin>:5043:12, :5054:12
      automatic logic [1:0][31:0] _T_82 = {{Register_inst80}, {_T_0}};	// <stdin>:5058:12, :5069:12
      automatic logic [1:0][31:0] _T_83 = {{Register_inst81}, {_T_0}};	// <stdin>:5073:12, :5084:12
      automatic logic [1:0][31:0] _T_84 = {{Register_inst82}, {_T_0}};	// <stdin>:5088:12, :5099:12
      automatic logic [1:0][31:0] _T_85 = {{Register_inst83}, {_T_0}};	// <stdin>:5103:12, :5114:12
      automatic logic [1:0][31:0] _T_86 = {{Register_inst84}, {_T_0}};	// <stdin>:5118:12, :5129:12
      automatic logic [1:0][31:0] _T_87 = {{Register_inst85}, {_T_0}};	// <stdin>:5133:12, :5144:12
      automatic logic [1:0][31:0] _T_88 = {{Register_inst86}, {_T_0}};	// <stdin>:5148:12, :5159:12
      automatic logic [1:0][31:0] _T_89 = {{Register_inst87}, {_T_0}};	// <stdin>:5163:12, :5174:12
      automatic logic [1:0][31:0] _T_90 = {{Register_inst88}, {_T_0}};	// <stdin>:5178:12, :5189:12
      automatic logic [1:0][31:0] _T_91 = {{Register_inst89}, {_T_0}};	// <stdin>:5193:12, :5204:12
      automatic logic [1:0][31:0] _T_92 = {{Register_inst90}, {_T_0}};	// <stdin>:5208:12, :5219:12
      automatic logic [1:0][31:0] _T_93 = {{Register_inst91}, {_T_0}};	// <stdin>:5223:12, :5234:12
      automatic logic [1:0][31:0] _T_94 = {{Register_inst92}, {_T_0}};	// <stdin>:5238:12, :5249:12
      automatic logic [1:0][31:0] _T_95 = {{Register_inst93}, {_T_0}};	// <stdin>:5253:12, :5264:12
      automatic logic [1:0][31:0] _T_96 = {{Register_inst94}, {_T_0}};	// <stdin>:5268:12, :5279:12
      automatic logic [1:0][31:0] _T_97 = {{Register_inst95}, {_T_0}};	// <stdin>:5283:12, :5294:12
      automatic logic [1:0][31:0] _T_98 = {{Register_inst96}, {_T_0}};	// <stdin>:5298:12, :5309:12
      automatic logic [1:0][31:0] _T_99 = {{Register_inst97}, {_T_0}};	// <stdin>:5313:12, :5324:12
      automatic logic [1:0][31:0] _T_100 = {{Register_inst98}, {_T_0}};	// <stdin>:5328:12, :5339:12
      automatic logic [1:0][31:0] _T_101 = {{Register_inst99}, {_T_0}};	// <stdin>:5343:12, :5354:12
      automatic logic [1:0][31:0] _T_102 = {{Register_inst100}, {_T_0}};	// <stdin>:5358:12, :5369:12
      automatic logic [1:0][31:0] _T_103 = {{Register_inst101}, {_T_0}};	// <stdin>:5373:12, :5384:12
      automatic logic [1:0][31:0] _T_104 = {{Register_inst102}, {_T_0}};	// <stdin>:5388:12, :5399:12
      automatic logic [1:0][31:0] _T_105 = {{Register_inst103}, {_T_0}};	// <stdin>:5403:12, :5414:12
      automatic logic [1:0][31:0] _T_106 = {{Register_inst104}, {_T_0}};	// <stdin>:5418:12, :5429:12
      automatic logic [1:0][31:0] _T_107 = {{Register_inst105}, {_T_0}};	// <stdin>:5433:12, :5444:12
      automatic logic [1:0][31:0] _T_108 = {{Register_inst106}, {_T_0}};	// <stdin>:5448:12, :5459:12
      automatic logic [1:0][31:0] _T_109 = {{Register_inst107}, {_T_0}};	// <stdin>:5463:12, :5474:12
      automatic logic [1:0][31:0] _T_110 = {{Register_inst108}, {_T_0}};	// <stdin>:5478:12, :5489:12
      automatic logic [1:0][31:0] _T_111 = {{Register_inst109}, {_T_0}};	// <stdin>:5493:12, :5504:12
      automatic logic [1:0][31:0] _T_112 = {{Register_inst110}, {_T_0}};	// <stdin>:5508:12, :5519:12
      automatic logic [1:0][31:0] _T_113 = {{Register_inst111}, {_T_0}};	// <stdin>:5523:12, :5534:12
      automatic logic [1:0][31:0] _T_114 = {{Register_inst112}, {_T_0}};	// <stdin>:5538:12, :5549:12
      automatic logic [1:0][31:0] _T_115 = {{Register_inst113}, {_T_0}};	// <stdin>:5553:12, :5564:12
      automatic logic [1:0][31:0] _T_116 = {{Register_inst114}, {_T_0}};	// <stdin>:5568:12, :5579:12
      automatic logic [1:0][31:0] _T_117 = {{Register_inst115}, {_T_0}};	// <stdin>:5583:12, :5594:12
      automatic logic [1:0][31:0] _T_118 = {{Register_inst116}, {_T_0}};	// <stdin>:5598:12, :5609:12
      automatic logic [1:0][31:0] _T_119 = {{Register_inst117}, {_T_0}};	// <stdin>:5613:12, :5624:12
      automatic logic [1:0][31:0] _T_120 = {{Register_inst118}, {_T_0}};	// <stdin>:5628:12, :5639:12
      automatic logic [1:0][31:0] _T_121 = {{Register_inst119}, {_T_0}};	// <stdin>:5643:12, :5654:12
      automatic logic [1:0][31:0] _T_122 = {{Register_inst120}, {_T_0}};	// <stdin>:5658:12, :5669:12
      automatic logic [1:0][31:0] _T_123 = {{Register_inst121}, {_T_0}};	// <stdin>:5673:12, :5684:12
      automatic logic [1:0][31:0] _T_124 = {{Register_inst122}, {_T_0}};	// <stdin>:5688:12, :5699:12
      automatic logic [1:0][31:0] _T_125 = {{Register_inst123}, {_T_0}};	// <stdin>:5703:12, :5714:12
      automatic logic [1:0][31:0] _T_126 = {{Register_inst124}, {_T_0}};	// <stdin>:5718:12, :5729:12
      automatic logic [1:0][31:0] _T_127 = {{Register_inst125}, {_T_0}};	// <stdin>:5733:12, :5744:12
      automatic logic [1:0][31:0] _T_128 = {{Register_inst126}, {_T_0}};	// <stdin>:5748:12, :5759:12
      automatic logic [1:0][31:0] _T_129 = {{Register_inst127}, {_T_0}};	// <stdin>:5763:12, :5774:12
      automatic logic [1:0][31:0] _T_130 = {{Register_inst128}, {_T_0}};	// <stdin>:5778:12, :5789:12
      automatic logic [1:0][31:0] _T_131 = {{Register_inst129}, {_T_0}};	// <stdin>:5793:12, :5804:12
      automatic logic [1:0][31:0] _T_132 = {{Register_inst130}, {_T_0}};	// <stdin>:5808:12, :5819:12
      automatic logic [1:0][31:0] _T_133 = {{Register_inst131}, {_T_0}};	// <stdin>:5823:12, :5834:12
      automatic logic [1:0][31:0] _T_134 = {{Register_inst132}, {_T_0}};	// <stdin>:5838:12, :5849:12
      automatic logic [1:0][31:0] _T_135 = {{Register_inst133}, {_T_0}};	// <stdin>:5853:12, :5864:12
      automatic logic [1:0][31:0] _T_136 = {{Register_inst134}, {_T_0}};	// <stdin>:5868:12, :5879:12
      automatic logic [1:0][31:0] _T_137 = {{Register_inst135}, {_T_0}};	// <stdin>:5883:12, :5894:12
      automatic logic [1:0][31:0] _T_138 = {{Register_inst136}, {_T_0}};	// <stdin>:5898:12, :5909:12
      automatic logic [1:0][31:0] _T_139 = {{Register_inst137}, {_T_0}};	// <stdin>:5913:12, :5924:12
      automatic logic [1:0][31:0] _T_140 = {{Register_inst138}, {_T_0}};	// <stdin>:5928:12, :5939:12
      automatic logic [1:0][31:0] _T_141 = {{Register_inst139}, {_T_0}};	// <stdin>:5943:12, :5954:12
      automatic logic [1:0][31:0] _T_142 = {{Register_inst140}, {_T_0}};	// <stdin>:5958:12, :5969:12
      automatic logic [1:0][31:0] _T_143 = {{Register_inst141}, {_T_0}};	// <stdin>:5973:12, :5984:12
      automatic logic [1:0][31:0] _T_144 = {{Register_inst142}, {_T_0}};	// <stdin>:5988:13, :5999:13
      automatic logic [1:0][31:0] _T_145 = {{Register_inst143}, {_T_0}};	// <stdin>:6003:13, :6014:13
      automatic logic [1:0][31:0] _T_146 = {{Register_inst144}, {_T_0}};	// <stdin>:6018:13, :6029:13
      automatic logic [1:0][31:0] _T_147 = {{Register_inst145}, {_T_0}};	// <stdin>:6033:13, :6044:13
      automatic logic [1:0][31:0] _T_148 = {{Register_inst146}, {_T_0}};	// <stdin>:6048:13, :6059:13
      automatic logic [1:0][31:0] _T_149 = {{Register_inst147}, {_T_0}};	// <stdin>:6063:13, :6074:13
      automatic logic [1:0][31:0] _T_150 = {{Register_inst148}, {_T_0}};	// <stdin>:6078:13, :6089:13
      automatic logic [1:0][31:0] _T_151 = {{Register_inst149}, {_T_0}};	// <stdin>:6093:13, :6104:13
      automatic logic [1:0][31:0] _T_152 = {{Register_inst150}, {_T_0}};	// <stdin>:6108:13, :6119:13
      automatic logic [1:0][31:0] _T_153 = {{Register_inst151}, {_T_0}};	// <stdin>:6123:13, :6134:13
      automatic logic [1:0][31:0] _T_154 = {{Register_inst152}, {_T_0}};	// <stdin>:6138:13, :6149:13
      automatic logic [1:0][31:0] _T_155 = {{Register_inst153}, {_T_0}};	// <stdin>:6153:13, :6164:13
      automatic logic [1:0][31:0] _T_156 = {{Register_inst154}, {_T_0}};	// <stdin>:6168:13, :6179:13
      automatic logic [1:0][31:0] _T_157 = {{Register_inst155}, {_T_0}};	// <stdin>:6183:13, :6194:13
      automatic logic [1:0][31:0] _T_158 = {{Register_inst156}, {_T_0}};	// <stdin>:6198:13, :6209:13
      automatic logic [1:0][31:0] _T_159 = {{Register_inst157}, {_T_0}};	// <stdin>:6213:13, :6224:13
      automatic logic [1:0][31:0] _T_160 = {{Register_inst158}, {_T_0}};	// <stdin>:6228:13, :6239:13
      automatic logic [1:0][31:0] _T_161 = {{Register_inst159}, {_T_0}};	// <stdin>:6243:13, :6254:13
      automatic logic [1:0][31:0] _T_162 = {{Register_inst160}, {_T_0}};	// <stdin>:6258:13, :6269:13
      automatic logic [1:0][31:0] _T_163 = {{Register_inst161}, {_T_0}};	// <stdin>:6273:13, :6284:13
      automatic logic [1:0][31:0] _T_164 = {{Register_inst162}, {_T_0}};	// <stdin>:6288:13, :6299:13
      automatic logic [1:0][31:0] _T_165 = {{Register_inst163}, {_T_0}};	// <stdin>:6303:13, :6314:13
      automatic logic [1:0][31:0] _T_166 = {{Register_inst164}, {_T_0}};	// <stdin>:6318:13, :6329:13
      automatic logic [1:0][31:0] _T_167 = {{Register_inst165}, {_T_0}};	// <stdin>:6333:13, :6344:13
      automatic logic [1:0][31:0] _T_168 = {{Register_inst166}, {_T_0}};	// <stdin>:6348:13, :6359:13
      automatic logic [1:0][31:0] _T_169 = {{Register_inst167}, {_T_0}};	// <stdin>:6363:13, :6374:13
      automatic logic [1:0][31:0] _T_170 = {{Register_inst168}, {_T_0}};	// <stdin>:6378:13, :6389:13
      automatic logic [1:0][31:0] _T_171 = {{Register_inst169}, {_T_0}};	// <stdin>:6393:13, :6404:13
      automatic logic [1:0][31:0] _T_172 = {{Register_inst170}, {_T_0}};	// <stdin>:6408:13, :6419:13
      automatic logic [1:0][31:0] _T_173 = {{Register_inst171}, {_T_0}};	// <stdin>:6423:13, :6434:13
      automatic logic [1:0][31:0] _T_174 = {{Register_inst172}, {_T_0}};	// <stdin>:6438:13, :6449:13
      automatic logic [1:0][31:0] _T_175 = {{Register_inst173}, {_T_0}};	// <stdin>:6453:13, :6464:13
      automatic logic [1:0][31:0] _T_176 = {{Register_inst174}, {_T_0}};	// <stdin>:6468:13, :6479:13
      automatic logic [1:0][31:0] _T_177 = {{Register_inst175}, {_T_0}};	// <stdin>:6483:13, :6494:13
      automatic logic [1:0][31:0] _T_178 = {{Register_inst176}, {_T_0}};	// <stdin>:6498:13, :6509:13
      automatic logic [1:0][31:0] _T_179 = {{Register_inst177}, {_T_0}};	// <stdin>:6513:13, :6524:13
      automatic logic [1:0][31:0] _T_180 = {{Register_inst178}, {_T_0}};	// <stdin>:6528:13, :6539:13
      automatic logic [1:0][31:0] _T_181 = {{Register_inst179}, {_T_0}};	// <stdin>:6543:13, :6554:13
      automatic logic [1:0][31:0] _T_182 = {{Register_inst180}, {_T_0}};	// <stdin>:6558:13, :6569:13
      automatic logic [1:0][31:0] _T_183 = {{Register_inst181}, {_T_0}};	// <stdin>:6573:13, :6584:13
      automatic logic [1:0][31:0] _T_184 = {{Register_inst182}, {_T_0}};	// <stdin>:6588:13, :6599:13
      automatic logic [1:0][31:0] _T_185 = {{Register_inst183}, {_T_0}};	// <stdin>:6603:13, :6614:13
      automatic logic [1:0][31:0] _T_186 = {{Register_inst184}, {_T_0}};	// <stdin>:6618:13, :6629:13
      automatic logic [1:0][31:0] _T_187 = {{Register_inst185}, {_T_0}};	// <stdin>:6633:13, :6644:13
      automatic logic [1:0][31:0] _T_188 = {{Register_inst186}, {_T_0}};	// <stdin>:6648:13, :6659:13
      automatic logic [1:0][31:0] _T_189 = {{Register_inst187}, {_T_0}};	// <stdin>:6663:13, :6674:13
      automatic logic [1:0][31:0] _T_190 = {{Register_inst188}, {_T_0}};	// <stdin>:6678:13, :6689:13
      automatic logic [1:0][31:0] _T_191 = {{Register_inst189}, {_T_0}};	// <stdin>:6693:13, :6704:13
      automatic logic [1:0][31:0] _T_192 = {{Register_inst190}, {_T_0}};	// <stdin>:6708:13, :6719:13
      automatic logic [1:0][31:0] _T_193 = {{Register_inst191}, {_T_0}};	// <stdin>:6723:13, :6734:13
      automatic logic [1:0][31:0] _T_194 = {{Register_inst192}, {_T_0}};	// <stdin>:6738:13, :6749:13
      automatic logic [1:0][31:0] _T_195 = {{Register_inst193}, {_T_0}};	// <stdin>:6753:13, :6764:13
      automatic logic [1:0][31:0] _T_196 = {{Register_inst194}, {_T_0}};	// <stdin>:6768:13, :6779:13
      automatic logic [1:0][31:0] _T_197 = {{Register_inst195}, {_T_0}};	// <stdin>:6783:13, :6794:13
      automatic logic [1:0][31:0] _T_198 = {{Register_inst196}, {_T_0}};	// <stdin>:6798:13, :6809:13
      automatic logic [1:0][31:0] _T_199 = {{Register_inst197}, {_T_0}};	// <stdin>:6813:13, :6824:13
      automatic logic [1:0][31:0] _T_200 = {{Register_inst198}, {_T_0}};	// <stdin>:6828:13, :6839:13
      automatic logic [1:0][31:0] _T_201 = {{Register_inst199}, {_T_0}};	// <stdin>:6843:13, :6854:13
      automatic logic [1:0][31:0] _T_202 = {{Register_inst200}, {_T_0}};	// <stdin>:6858:13, :6869:13
      automatic logic [1:0][31:0] _T_203 = {{Register_inst201}, {_T_0}};	// <stdin>:6873:13, :6884:13
      automatic logic [1:0][31:0] _T_204 = {{Register_inst202}, {_T_0}};	// <stdin>:6888:13, :6899:13
      automatic logic [1:0][31:0] _T_205 = {{Register_inst203}, {_T_0}};	// <stdin>:6903:13, :6914:13
      automatic logic [1:0][31:0] _T_206 = {{Register_inst204}, {_T_0}};	// <stdin>:6918:13, :6929:13
      automatic logic [1:0][31:0] _T_207 = {{Register_inst205}, {_T_0}};	// <stdin>:6933:13, :6944:13
      automatic logic [1:0][31:0] _T_208 = {{Register_inst206}, {_T_0}};	// <stdin>:6948:13, :6959:13
      automatic logic [1:0][31:0] _T_209 = {{Register_inst207}, {_T_0}};	// <stdin>:6963:13, :6974:13
      automatic logic [1:0][31:0] _T_210 = {{Register_inst208}, {_T_0}};	// <stdin>:6978:13, :6989:13
      automatic logic [1:0][31:0] _T_211 = {{Register_inst209}, {_T_0}};	// <stdin>:6993:13, :7004:13
      automatic logic [1:0][31:0] _T_212 = {{Register_inst210}, {_T_0}};	// <stdin>:7008:13, :7019:13
      automatic logic [1:0][31:0] _T_213 = {{Register_inst211}, {_T_0}};	// <stdin>:7023:13, :7034:13
      automatic logic [1:0][31:0] _T_214 = {{Register_inst212}, {_T_0}};	// <stdin>:7038:13, :7049:13
      automatic logic [1:0][31:0] _T_215 = {{Register_inst213}, {_T_0}};	// <stdin>:7053:13, :7064:13
      automatic logic [1:0][31:0] _T_216 = {{Register_inst214}, {_T_0}};	// <stdin>:7068:13, :7079:13
      automatic logic [1:0][31:0] _T_217 = {{Register_inst215}, {_T_0}};	// <stdin>:7083:13, :7094:13
      automatic logic [1:0][31:0] _T_218 = {{Register_inst216}, {_T_0}};	// <stdin>:7098:13, :7109:13
      automatic logic [1:0][31:0] _T_219 = {{Register_inst217}, {_T_0}};	// <stdin>:7113:13, :7124:13
      automatic logic [1:0][31:0] _T_220 = {{Register_inst218}, {_T_0}};	// <stdin>:7128:13, :7139:13
      automatic logic [1:0][31:0] _T_221 = {{Register_inst219}, {_T_0}};	// <stdin>:7143:13, :7154:13
      automatic logic [1:0][31:0] _T_222 = {{Register_inst220}, {_T_0}};	// <stdin>:7158:13, :7169:13
      automatic logic [1:0][31:0] _T_223 = {{Register_inst221}, {_T_0}};	// <stdin>:7173:13, :7184:13
      automatic logic [1:0][31:0] _T_224 = {{Register_inst222}, {_T_0}};	// <stdin>:7188:13, :7199:13
      automatic logic [1:0][31:0] _T_225 = {{Register_inst223}, {_T_0}};	// <stdin>:7203:13, :7214:13
      automatic logic [1:0][31:0] _T_226 = {{Register_inst224}, {_T_0}};	// <stdin>:7218:13, :7229:13
      automatic logic [1:0][31:0] _T_227 = {{Register_inst225}, {_T_0}};	// <stdin>:7233:13, :7244:13
      automatic logic [1:0][31:0] _T_228 = {{Register_inst226}, {_T_0}};	// <stdin>:7248:13, :7259:13
      automatic logic [1:0][31:0] _T_229 = {{Register_inst227}, {_T_0}};	// <stdin>:7263:13, :7274:13
      automatic logic [1:0][31:0] _T_230 = {{Register_inst228}, {_T_0}};	// <stdin>:7278:13, :7289:13
      automatic logic [1:0][31:0] _T_231 = {{Register_inst229}, {_T_0}};	// <stdin>:7293:13, :7304:13
      automatic logic [1:0][31:0] _T_232 = {{Register_inst230}, {_T_0}};	// <stdin>:7308:13, :7319:13
      automatic logic [1:0][31:0] _T_233 = {{Register_inst231}, {_T_0}};	// <stdin>:7323:13, :7334:13
      automatic logic [1:0][31:0] _T_234 = {{Register_inst232}, {_T_0}};	// <stdin>:7338:13, :7349:13
      automatic logic [1:0][31:0] _T_235 = {{Register_inst233}, {_T_0}};	// <stdin>:7353:13, :7364:13
      automatic logic [1:0][31:0] _T_236 = {{Register_inst234}, {_T_0}};	// <stdin>:7368:13, :7379:13
      automatic logic [1:0][31:0] _T_237 = {{Register_inst235}, {_T_0}};	// <stdin>:7383:13, :7394:13
      automatic logic [1:0][31:0] _T_238 = {{Register_inst236}, {_T_0}};	// <stdin>:7398:13, :7409:13
      automatic logic [1:0][31:0] _T_239 = {{Register_inst237}, {_T_0}};	// <stdin>:7413:13, :7424:13
      automatic logic [1:0][31:0] _T_240 = {{Register_inst238}, {_T_0}};	// <stdin>:7428:13, :7439:13
      automatic logic [1:0][31:0] _T_241 = {{Register_inst239}, {_T_0}};	// <stdin>:7443:13, :7454:13
      automatic logic [1:0][31:0] _T_242 = {{Register_inst240}, {_T_0}};	// <stdin>:7458:13, :7469:13
      automatic logic [1:0][31:0] _T_243 = {{Register_inst241}, {_T_0}};	// <stdin>:7473:13, :7484:13
      automatic logic [1:0][31:0] _T_244 = {{Register_inst242}, {_T_0}};	// <stdin>:7488:13, :7499:13
      automatic logic [1:0][31:0] _T_245 = {{Register_inst243}, {_T_0}};	// <stdin>:7503:13, :7514:13
      automatic logic [1:0][31:0] _T_246 = {{Register_inst244}, {_T_0}};	// <stdin>:7518:13, :7529:13
      automatic logic [1:0][31:0] _T_247 = {{Register_inst245}, {_T_0}};	// <stdin>:7533:13, :7544:13
      automatic logic [1:0][31:0] _T_248 = {{Register_inst246}, {_T_0}};	// <stdin>:7548:13, :7559:13
      automatic logic [1:0][31:0] _T_249 = {{Register_inst247}, {_T_0}};	// <stdin>:7563:13, :7574:13
      automatic logic [1:0][31:0] _T_250 = {{Register_inst248}, {_T_0}};	// <stdin>:7578:13, :7589:13
      automatic logic [1:0][31:0] _T_251 = {{Register_inst249}, {_T_0}};	// <stdin>:7593:13, :7604:13
      automatic logic [1:0][31:0] _T_252 = {{Register_inst250}, {_T_0}};	// <stdin>:7608:13, :7619:13
      automatic logic [1:0][31:0] _T_253 = {{Register_inst251}, {_T_0}};	// <stdin>:7623:13, :7634:13
      automatic logic [1:0][31:0] _T_254 = {{Register_inst252}, {_T_0}};	// <stdin>:7638:13, :7649:13
      automatic logic [1:0][31:0] _T_255 = {{Register_inst253}, {_T_0}};	// <stdin>:7653:13, :7664:13
      automatic logic [1:0][31:0] _T_256 = {{Register_inst254}, {_T_0}};	// <stdin>:7668:13, :7679:13
      automatic logic [1:0][31:0] _T_257 = {{Register_inst255}, {_T_0}};	// <stdin>:7683:13, :7694:13

      Register_inst0 <= _T_2[_T_1 == 8'h0 & write_0_en];	// <stdin>:3854:10, :3855:10, :3856:10, :3858:10, :3861:9
      Register_inst1 <= _T_3[_T_1 == 8'h1 & write_0_en];	// <stdin>:3870:11, :3871:11, :3872:11, :3874:11, :3877:9
      Register_inst2 <= _T_4[_T_1 == 8'h2 & write_0_en];	// <stdin>:3885:11, :3886:11, :3887:11, :3889:11, :3892:9
      Register_inst3 <= _T_5[_T_1 == 8'h3 & write_0_en];	// <stdin>:3900:11, :3901:11, :3902:11, :3904:11, :3907:9
      Register_inst4 <= _T_6[_T_1 == 8'h4 & write_0_en];	// <stdin>:3915:11, :3916:11, :3917:11, :3919:11, :3922:9
      Register_inst5 <= _T_7[_T_1 == 8'h5 & write_0_en];	// <stdin>:3930:11, :3931:11, :3932:11, :3934:11, :3937:9
      Register_inst6 <= _T_8[_T_1 == 8'h6 & write_0_en];	// <stdin>:3945:11, :3946:11, :3947:11, :3949:11, :3952:9
      Register_inst7 <= _T_9[_T_1 == 8'h7 & write_0_en];	// <stdin>:3960:11, :3961:11, :3962:11, :3964:11, :3967:9
      Register_inst8 <= _T_10[_T_1 == 8'h8 & write_0_en];	// <stdin>:3975:11, :3976:11, :3977:11, :3979:11, :3982:9
      Register_inst9 <= _T_11[_T_1 == 8'h9 & write_0_en];	// <stdin>:3990:11, :3991:11, :3992:11, :3994:11, :3997:9
      Register_inst10 <= _T_12[_T_1 == 8'hA & write_0_en];	// <stdin>:4005:11, :4006:11, :4007:11, :4009:11, :4012:9
      Register_inst11 <= _T_13[_T_1 == 8'hB & write_0_en];	// <stdin>:4020:11, :4021:11, :4022:11, :4024:11, :4027:9
      Register_inst12 <= _T_14[_T_1 == 8'hC & write_0_en];	// <stdin>:4035:11, :4036:11, :4037:11, :4039:11, :4042:9
      Register_inst13 <= _T_15[_T_1 == 8'hD & write_0_en];	// <stdin>:4050:11, :4051:11, :4052:11, :4054:11, :4057:9
      Register_inst14 <= _T_16[_T_1 == 8'hE & write_0_en];	// <stdin>:4065:12, :4066:12, :4067:12, :4069:12, :4072:9
      Register_inst15 <= _T_17[_T_1 == 8'hF & write_0_en];	// <stdin>:4080:12, :4081:12, :4082:12, :4084:12, :4087:9
      Register_inst16 <= _T_18[_T_1 == 8'h10 & write_0_en];	// <stdin>:4095:12, :4096:12, :4097:12, :4099:12, :4102:9
      Register_inst17 <= _T_19[_T_1 == 8'h11 & write_0_en];	// <stdin>:4110:12, :4111:12, :4112:12, :4114:12, :4117:9
      Register_inst18 <= _T_20[_T_1 == 8'h12 & write_0_en];	// <stdin>:4125:12, :4126:12, :4127:12, :4129:12, :4132:9
      Register_inst19 <= _T_21[_T_1 == 8'h13 & write_0_en];	// <stdin>:4140:12, :4141:12, :4142:12, :4144:12, :4147:9
      Register_inst20 <= _T_22[_T_1 == 8'h14 & write_0_en];	// <stdin>:4155:12, :4156:12, :4157:12, :4159:12, :4162:9
      Register_inst21 <= _T_23[_T_1 == 8'h15 & write_0_en];	// <stdin>:4170:12, :4171:12, :4172:12, :4174:12, :4177:9
      Register_inst22 <= _T_24[_T_1 == 8'h16 & write_0_en];	// <stdin>:4185:12, :4186:12, :4187:12, :4189:12, :4192:9
      Register_inst23 <= _T_25[_T_1 == 8'h17 & write_0_en];	// <stdin>:4200:12, :4201:12, :4202:12, :4204:12, :4207:9
      Register_inst24 <= _T_26[_T_1 == 8'h18 & write_0_en];	// <stdin>:4215:12, :4216:12, :4217:12, :4219:12, :4222:9
      Register_inst25 <= _T_27[_T_1 == 8'h19 & write_0_en];	// <stdin>:4230:12, :4231:12, :4232:12, :4234:12, :4237:9
      Register_inst26 <= _T_28[_T_1 == 8'h1A & write_0_en];	// <stdin>:4245:12, :4246:12, :4247:12, :4249:12, :4252:9
      Register_inst27 <= _T_29[_T_1 == 8'h1B & write_0_en];	// <stdin>:4260:12, :4261:12, :4262:12, :4264:12, :4267:9
      Register_inst28 <= _T_30[_T_1 == 8'h1C & write_0_en];	// <stdin>:4275:12, :4276:12, :4277:12, :4279:12, :4282:9
      Register_inst29 <= _T_31[_T_1 == 8'h1D & write_0_en];	// <stdin>:4290:12, :4291:12, :4292:12, :4294:12, :4297:9
      Register_inst30 <= _T_32[_T_1 == 8'h1E & write_0_en];	// <stdin>:4305:12, :4306:12, :4307:12, :4309:12, :4312:9
      Register_inst31 <= _T_33[_T_1 == 8'h1F & write_0_en];	// <stdin>:4320:12, :4321:12, :4322:12, :4324:12, :4327:9
      Register_inst32 <= _T_34[_T_1 == 8'h20 & write_0_en];	// <stdin>:4335:12, :4336:12, :4337:12, :4339:12, :4342:9
      Register_inst33 <= _T_35[_T_1 == 8'h21 & write_0_en];	// <stdin>:4350:12, :4351:12, :4352:12, :4354:12, :4357:9
      Register_inst34 <= _T_36[_T_1 == 8'h22 & write_0_en];	// <stdin>:4365:12, :4366:12, :4367:12, :4369:12, :4372:9
      Register_inst35 <= _T_37[_T_1 == 8'h23 & write_0_en];	// <stdin>:4380:12, :4381:12, :4382:12, :4384:12, :4387:9
      Register_inst36 <= _T_38[_T_1 == 8'h24 & write_0_en];	// <stdin>:4395:12, :4396:12, :4397:12, :4399:12, :4402:9
      Register_inst37 <= _T_39[_T_1 == 8'h25 & write_0_en];	// <stdin>:4410:12, :4411:12, :4412:12, :4414:12, :4417:9
      Register_inst38 <= _T_40[_T_1 == 8'h26 & write_0_en];	// <stdin>:4425:12, :4426:12, :4427:12, :4429:12, :4432:9
      Register_inst39 <= _T_41[_T_1 == 8'h27 & write_0_en];	// <stdin>:4440:12, :4441:12, :4442:12, :4444:12, :4447:9
      Register_inst40 <= _T_42[_T_1 == 8'h28 & write_0_en];	// <stdin>:4455:12, :4456:12, :4457:12, :4459:12, :4462:9
      Register_inst41 <= _T_43[_T_1 == 8'h29 & write_0_en];	// <stdin>:4470:12, :4471:12, :4472:12, :4474:12, :4477:9
      Register_inst42 <= _T_44[_T_1 == 8'h2A & write_0_en];	// <stdin>:4485:12, :4486:12, :4487:12, :4489:12, :4492:9
      Register_inst43 <= _T_45[_T_1 == 8'h2B & write_0_en];	// <stdin>:4500:12, :4501:12, :4502:12, :4504:12, :4507:9
      Register_inst44 <= _T_46[_T_1 == 8'h2C & write_0_en];	// <stdin>:4515:12, :4516:12, :4517:12, :4519:12, :4522:9
      Register_inst45 <= _T_47[_T_1 == 8'h2D & write_0_en];	// <stdin>:4530:12, :4531:12, :4532:12, :4534:12, :4537:9
      Register_inst46 <= _T_48[_T_1 == 8'h2E & write_0_en];	// <stdin>:4545:12, :4546:12, :4547:12, :4549:12, :4552:9
      Register_inst47 <= _T_49[_T_1 == 8'h2F & write_0_en];	// <stdin>:4560:12, :4561:12, :4562:12, :4564:12, :4567:9
      Register_inst48 <= _T_50[_T_1 == 8'h30 & write_0_en];	// <stdin>:4575:12, :4576:12, :4577:12, :4579:12, :4582:9
      Register_inst49 <= _T_51[_T_1 == 8'h31 & write_0_en];	// <stdin>:4590:12, :4591:12, :4592:12, :4594:12, :4597:9
      Register_inst50 <= _T_52[_T_1 == 8'h32 & write_0_en];	// <stdin>:4605:12, :4606:12, :4607:12, :4609:12, :4612:9
      Register_inst51 <= _T_53[_T_1 == 8'h33 & write_0_en];	// <stdin>:4620:12, :4621:12, :4622:12, :4624:12, :4627:9
      Register_inst52 <= _T_54[_T_1 == 8'h34 & write_0_en];	// <stdin>:4635:12, :4636:12, :4637:12, :4639:12, :4642:9
      Register_inst53 <= _T_55[_T_1 == 8'h35 & write_0_en];	// <stdin>:4650:12, :4651:12, :4652:12, :4654:12, :4657:9
      Register_inst54 <= _T_56[_T_1 == 8'h36 & write_0_en];	// <stdin>:4665:12, :4666:12, :4667:12, :4669:12, :4672:9
      Register_inst55 <= _T_57[_T_1 == 8'h37 & write_0_en];	// <stdin>:4680:12, :4681:12, :4682:12, :4684:12, :4687:9
      Register_inst56 <= _T_58[_T_1 == 8'h38 & write_0_en];	// <stdin>:4695:12, :4696:12, :4697:12, :4699:12, :4702:9
      Register_inst57 <= _T_59[_T_1 == 8'h39 & write_0_en];	// <stdin>:4710:12, :4711:12, :4712:12, :4714:12, :4717:9
      Register_inst58 <= _T_60[_T_1 == 8'h3A & write_0_en];	// <stdin>:4725:12, :4726:12, :4727:12, :4729:12, :4732:9
      Register_inst59 <= _T_61[_T_1 == 8'h3B & write_0_en];	// <stdin>:4740:12, :4741:12, :4742:12, :4744:12, :4747:9
      Register_inst60 <= _T_62[_T_1 == 8'h3C & write_0_en];	// <stdin>:4755:12, :4756:12, :4757:12, :4759:12, :4762:9
      Register_inst61 <= _T_63[_T_1 == 8'h3D & write_0_en];	// <stdin>:4770:12, :4771:12, :4772:12, :4774:12, :4777:9
      Register_inst62 <= _T_64[_T_1 == 8'h3E & write_0_en];	// <stdin>:4785:12, :4786:12, :4787:12, :4789:12, :4792:9
      Register_inst63 <= _T_65[_T_1 == 8'h3F & write_0_en];	// <stdin>:4800:12, :4801:12, :4802:12, :4804:12, :4807:9
      Register_inst64 <= _T_66[_T_1 == 8'h40 & write_0_en];	// <stdin>:4815:12, :4816:12, :4817:12, :4819:12, :4822:9
      Register_inst65 <= _T_67[_T_1 == 8'h41 & write_0_en];	// <stdin>:4830:12, :4831:12, :4832:12, :4834:12, :4837:9
      Register_inst66 <= _T_68[_T_1 == 8'h42 & write_0_en];	// <stdin>:4845:12, :4846:12, :4847:12, :4849:12, :4852:9
      Register_inst67 <= _T_69[_T_1 == 8'h43 & write_0_en];	// <stdin>:4860:12, :4861:12, :4862:12, :4864:12, :4867:9
      Register_inst68 <= _T_70[_T_1 == 8'h44 & write_0_en];	// <stdin>:4875:12, :4876:12, :4877:12, :4879:12, :4882:9
      Register_inst69 <= _T_71[_T_1 == 8'h45 & write_0_en];	// <stdin>:4890:12, :4891:12, :4892:12, :4894:12, :4897:9
      Register_inst70 <= _T_72[_T_1 == 8'h46 & write_0_en];	// <stdin>:4905:12, :4906:12, :4907:12, :4909:12, :4912:9
      Register_inst71 <= _T_73[_T_1 == 8'h47 & write_0_en];	// <stdin>:4920:12, :4921:12, :4922:12, :4924:12, :4927:9
      Register_inst72 <= _T_74[_T_1 == 8'h48 & write_0_en];	// <stdin>:4935:12, :4936:12, :4937:12, :4939:12, :4942:9
      Register_inst73 <= _T_75[_T_1 == 8'h49 & write_0_en];	// <stdin>:4950:12, :4951:12, :4952:12, :4954:12, :4957:9
      Register_inst74 <= _T_76[_T_1 == 8'h4A & write_0_en];	// <stdin>:4965:12, :4966:12, :4967:12, :4969:12, :4972:9
      Register_inst75 <= _T_77[_T_1 == 8'h4B & write_0_en];	// <stdin>:4980:12, :4981:12, :4982:12, :4984:12, :4987:9
      Register_inst76 <= _T_78[_T_1 == 8'h4C & write_0_en];	// <stdin>:4995:12, :4996:12, :4997:12, :4999:12, :5002:9
      Register_inst77 <= _T_79[_T_1 == 8'h4D & write_0_en];	// <stdin>:5010:12, :5011:12, :5012:12, :5014:12, :5017:9
      Register_inst78 <= _T_80[_T_1 == 8'h4E & write_0_en];	// <stdin>:5025:12, :5026:12, :5027:12, :5029:12, :5032:9
      Register_inst79 <= _T_81[_T_1 == 8'h4F & write_0_en];	// <stdin>:5040:12, :5041:12, :5042:12, :5044:12, :5047:9
      Register_inst80 <= _T_82[_T_1 == 8'h50 & write_0_en];	// <stdin>:5055:12, :5056:12, :5057:12, :5059:12, :5062:9
      Register_inst81 <= _T_83[_T_1 == 8'h51 & write_0_en];	// <stdin>:5070:12, :5071:12, :5072:12, :5074:12, :5077:9
      Register_inst82 <= _T_84[_T_1 == 8'h52 & write_0_en];	// <stdin>:5085:12, :5086:12, :5087:12, :5089:12, :5092:9
      Register_inst83 <= _T_85[_T_1 == 8'h53 & write_0_en];	// <stdin>:5100:12, :5101:12, :5102:12, :5104:12, :5107:9
      Register_inst84 <= _T_86[_T_1 == 8'h54 & write_0_en];	// <stdin>:5115:12, :5116:12, :5117:12, :5119:12, :5122:9
      Register_inst85 <= _T_87[_T_1 == 8'h55 & write_0_en];	// <stdin>:5130:12, :5131:12, :5132:12, :5134:12, :5137:9
      Register_inst86 <= _T_88[_T_1 == 8'h56 & write_0_en];	// <stdin>:5145:12, :5146:12, :5147:12, :5149:12, :5152:9
      Register_inst87 <= _T_89[_T_1 == 8'h57 & write_0_en];	// <stdin>:5160:12, :5161:12, :5162:12, :5164:12, :5167:9
      Register_inst88 <= _T_90[_T_1 == 8'h58 & write_0_en];	// <stdin>:5175:12, :5176:12, :5177:12, :5179:12, :5182:9
      Register_inst89 <= _T_91[_T_1 == 8'h59 & write_0_en];	// <stdin>:5190:12, :5191:12, :5192:12, :5194:12, :5197:9
      Register_inst90 <= _T_92[_T_1 == 8'h5A & write_0_en];	// <stdin>:5205:12, :5206:12, :5207:12, :5209:12, :5212:9
      Register_inst91 <= _T_93[_T_1 == 8'h5B & write_0_en];	// <stdin>:5220:12, :5221:12, :5222:12, :5224:12, :5227:9
      Register_inst92 <= _T_94[_T_1 == 8'h5C & write_0_en];	// <stdin>:5235:12, :5236:12, :5237:12, :5239:12, :5242:9
      Register_inst93 <= _T_95[_T_1 == 8'h5D & write_0_en];	// <stdin>:5250:12, :5251:12, :5252:12, :5254:12, :5257:9
      Register_inst94 <= _T_96[_T_1 == 8'h5E & write_0_en];	// <stdin>:5265:12, :5266:12, :5267:12, :5269:12, :5272:9
      Register_inst95 <= _T_97[_T_1 == 8'h5F & write_0_en];	// <stdin>:5280:12, :5281:12, :5282:12, :5284:12, :5287:9
      Register_inst96 <= _T_98[_T_1 == 8'h60 & write_0_en];	// <stdin>:5295:12, :5296:12, :5297:12, :5299:12, :5302:9
      Register_inst97 <= _T_99[_T_1 == 8'h61 & write_0_en];	// <stdin>:5310:12, :5311:12, :5312:12, :5314:12, :5317:9
      Register_inst98 <= _T_100[_T_1 == 8'h62 & write_0_en];	// <stdin>:5325:12, :5326:12, :5327:12, :5329:12, :5332:9
      Register_inst99 <= _T_101[_T_1 == 8'h63 & write_0_en];	// <stdin>:5340:12, :5341:12, :5342:12, :5344:12, :5347:9
      Register_inst100 <= _T_102[_T_1 == 8'h64 & write_0_en];	// <stdin>:5355:12, :5356:12, :5357:12, :5359:12, :5362:9
      Register_inst101 <= _T_103[_T_1 == 8'h65 & write_0_en];	// <stdin>:5370:12, :5371:12, :5372:12, :5374:12, :5377:9
      Register_inst102 <= _T_104[_T_1 == 8'h66 & write_0_en];	// <stdin>:5385:12, :5386:12, :5387:12, :5389:12, :5392:9
      Register_inst103 <= _T_105[_T_1 == 8'h67 & write_0_en];	// <stdin>:5400:12, :5401:12, :5402:12, :5404:12, :5407:9
      Register_inst104 <= _T_106[_T_1 == 8'h68 & write_0_en];	// <stdin>:5415:12, :5416:12, :5417:12, :5419:12, :5422:9
      Register_inst105 <= _T_107[_T_1 == 8'h69 & write_0_en];	// <stdin>:5430:12, :5431:12, :5432:12, :5434:12, :5437:9
      Register_inst106 <= _T_108[_T_1 == 8'h6A & write_0_en];	// <stdin>:5445:12, :5446:12, :5447:12, :5449:12, :5452:9
      Register_inst107 <= _T_109[_T_1 == 8'h6B & write_0_en];	// <stdin>:5460:12, :5461:12, :5462:12, :5464:12, :5467:9
      Register_inst108 <= _T_110[_T_1 == 8'h6C & write_0_en];	// <stdin>:5475:12, :5476:12, :5477:12, :5479:12, :5482:9
      Register_inst109 <= _T_111[_T_1 == 8'h6D & write_0_en];	// <stdin>:5490:12, :5491:12, :5492:12, :5494:12, :5497:9
      Register_inst110 <= _T_112[_T_1 == 8'h6E & write_0_en];	// <stdin>:5505:12, :5506:12, :5507:12, :5509:12, :5512:9
      Register_inst111 <= _T_113[_T_1 == 8'h6F & write_0_en];	// <stdin>:5520:12, :5521:12, :5522:12, :5524:12, :5527:9
      Register_inst112 <= _T_114[_T_1 == 8'h70 & write_0_en];	// <stdin>:5535:12, :5536:12, :5537:12, :5539:12, :5542:9
      Register_inst113 <= _T_115[_T_1 == 8'h71 & write_0_en];	// <stdin>:5550:12, :5551:12, :5552:12, :5554:12, :5557:9
      Register_inst114 <= _T_116[_T_1 == 8'h72 & write_0_en];	// <stdin>:5565:12, :5566:12, :5567:12, :5569:12, :5572:9
      Register_inst115 <= _T_117[_T_1 == 8'h73 & write_0_en];	// <stdin>:5580:12, :5581:12, :5582:12, :5584:12, :5587:9
      Register_inst116 <= _T_118[_T_1 == 8'h74 & write_0_en];	// <stdin>:5595:12, :5596:12, :5597:12, :5599:12, :5602:9
      Register_inst117 <= _T_119[_T_1 == 8'h75 & write_0_en];	// <stdin>:5610:12, :5611:12, :5612:12, :5614:12, :5617:9
      Register_inst118 <= _T_120[_T_1 == 8'h76 & write_0_en];	// <stdin>:5625:12, :5626:12, :5627:12, :5629:12, :5632:9
      Register_inst119 <= _T_121[_T_1 == 8'h77 & write_0_en];	// <stdin>:5640:12, :5641:12, :5642:12, :5644:12, :5647:9
      Register_inst120 <= _T_122[_T_1 == 8'h78 & write_0_en];	// <stdin>:5655:12, :5656:12, :5657:12, :5659:12, :5662:9
      Register_inst121 <= _T_123[_T_1 == 8'h79 & write_0_en];	// <stdin>:5670:12, :5671:12, :5672:12, :5674:12, :5677:9
      Register_inst122 <= _T_124[_T_1 == 8'h7A & write_0_en];	// <stdin>:5685:12, :5686:12, :5687:12, :5689:12, :5692:9
      Register_inst123 <= _T_125[_T_1 == 8'h7B & write_0_en];	// <stdin>:5700:12, :5701:12, :5702:12, :5704:12, :5707:9
      Register_inst124 <= _T_126[_T_1 == 8'h7C & write_0_en];	// <stdin>:5715:12, :5716:12, :5717:12, :5719:12, :5722:9
      Register_inst125 <= _T_127[_T_1 == 8'h7D & write_0_en];	// <stdin>:5730:12, :5731:12, :5732:12, :5734:12, :5737:9
      Register_inst126 <= _T_128[_T_1 == 8'h7E & write_0_en];	// <stdin>:5745:12, :5746:12, :5747:12, :5749:12, :5752:9
      Register_inst127 <= _T_129[_T_1 == 8'h7F & write_0_en];	// <stdin>:5760:12, :5761:12, :5762:12, :5764:12, :5767:9
      Register_inst128 <= _T_130[_T_1 == 8'h80 & write_0_en];	// <stdin>:5775:12, :5776:12, :5777:12, :5779:12, :5782:9
      Register_inst129 <= _T_131[_T_1 == 8'h81 & write_0_en];	// <stdin>:5790:12, :5791:12, :5792:12, :5794:12, :5797:9
      Register_inst130 <= _T_132[_T_1 == 8'h82 & write_0_en];	// <stdin>:5805:12, :5806:12, :5807:12, :5809:12, :5812:9
      Register_inst131 <= _T_133[_T_1 == 8'h83 & write_0_en];	// <stdin>:5820:12, :5821:12, :5822:12, :5824:12, :5827:9
      Register_inst132 <= _T_134[_T_1 == 8'h84 & write_0_en];	// <stdin>:5835:12, :5836:12, :5837:12, :5839:12, :5842:9
      Register_inst133 <= _T_135[_T_1 == 8'h85 & write_0_en];	// <stdin>:5850:12, :5851:12, :5852:12, :5854:12, :5857:9
      Register_inst134 <= _T_136[_T_1 == 8'h86 & write_0_en];	// <stdin>:5865:12, :5866:12, :5867:12, :5869:12, :5872:9
      Register_inst135 <= _T_137[_T_1 == 8'h87 & write_0_en];	// <stdin>:5880:12, :5881:12, :5882:12, :5884:12, :5887:9
      Register_inst136 <= _T_138[_T_1 == 8'h88 & write_0_en];	// <stdin>:5895:12, :5896:12, :5897:12, :5899:12, :5902:9
      Register_inst137 <= _T_139[_T_1 == 8'h89 & write_0_en];	// <stdin>:5910:12, :5911:12, :5912:12, :5914:12, :5917:9
      Register_inst138 <= _T_140[_T_1 == 8'h8A & write_0_en];	// <stdin>:5925:12, :5926:12, :5927:12, :5929:12, :5932:9
      Register_inst139 <= _T_141[_T_1 == 8'h8B & write_0_en];	// <stdin>:5940:12, :5941:12, :5942:12, :5944:12, :5947:9
      Register_inst140 <= _T_142[_T_1 == 8'h8C & write_0_en];	// <stdin>:5955:12, :5956:12, :5957:12, :5959:12, :5962:9
      Register_inst141 <= _T_143[_T_1 == 8'h8D & write_0_en];	// <stdin>:5970:12, :5971:12, :5972:12, :5974:12, :5977:9
      Register_inst142 <= _T_144[_T_1 == 8'h8E & write_0_en];	// <stdin>:5985:12, :5986:12, :5987:12, :5989:13, :5992:9
      Register_inst143 <= _T_145[_T_1 == 8'h8F & write_0_en];	// <stdin>:6000:13, :6001:13, :6002:13, :6004:13, :6007:9
      Register_inst144 <= _T_146[_T_1 == 8'h90 & write_0_en];	// <stdin>:6015:13, :6016:13, :6017:13, :6019:13, :6022:9
      Register_inst145 <= _T_147[_T_1 == 8'h91 & write_0_en];	// <stdin>:6030:13, :6031:13, :6032:13, :6034:13, :6037:9
      Register_inst146 <= _T_148[_T_1 == 8'h92 & write_0_en];	// <stdin>:6045:13, :6046:13, :6047:13, :6049:13, :6052:9
      Register_inst147 <= _T_149[_T_1 == 8'h93 & write_0_en];	// <stdin>:6060:13, :6061:13, :6062:13, :6064:13, :6067:9
      Register_inst148 <= _T_150[_T_1 == 8'h94 & write_0_en];	// <stdin>:6075:13, :6076:13, :6077:13, :6079:13, :6082:9
      Register_inst149 <= _T_151[_T_1 == 8'h95 & write_0_en];	// <stdin>:6090:13, :6091:13, :6092:13, :6094:13, :6097:9
      Register_inst150 <= _T_152[_T_1 == 8'h96 & write_0_en];	// <stdin>:6105:13, :6106:13, :6107:13, :6109:13, :6112:9
      Register_inst151 <= _T_153[_T_1 == 8'h97 & write_0_en];	// <stdin>:6120:13, :6121:13, :6122:13, :6124:13, :6127:9
      Register_inst152 <= _T_154[_T_1 == 8'h98 & write_0_en];	// <stdin>:6135:13, :6136:13, :6137:13, :6139:13, :6142:9
      Register_inst153 <= _T_155[_T_1 == 8'h99 & write_0_en];	// <stdin>:6150:13, :6151:13, :6152:13, :6154:13, :6157:9
      Register_inst154 <= _T_156[_T_1 == 8'h9A & write_0_en];	// <stdin>:6165:13, :6166:13, :6167:13, :6169:13, :6172:9
      Register_inst155 <= _T_157[_T_1 == 8'h9B & write_0_en];	// <stdin>:6180:13, :6181:13, :6182:13, :6184:13, :6187:9
      Register_inst156 <= _T_158[_T_1 == 8'h9C & write_0_en];	// <stdin>:6195:13, :6196:13, :6197:13, :6199:13, :6202:9
      Register_inst157 <= _T_159[_T_1 == 8'h9D & write_0_en];	// <stdin>:6210:13, :6211:13, :6212:13, :6214:13, :6217:9
      Register_inst158 <= _T_160[_T_1 == 8'h9E & write_0_en];	// <stdin>:6225:13, :6226:13, :6227:13, :6229:13, :6232:9
      Register_inst159 <= _T_161[_T_1 == 8'h9F & write_0_en];	// <stdin>:6240:13, :6241:13, :6242:13, :6244:13, :6247:9
      Register_inst160 <= _T_162[_T_1 == 8'hA0 & write_0_en];	// <stdin>:6255:13, :6256:13, :6257:13, :6259:13, :6262:9
      Register_inst161 <= _T_163[_T_1 == 8'hA1 & write_0_en];	// <stdin>:6270:13, :6271:13, :6272:13, :6274:13, :6277:9
      Register_inst162 <= _T_164[_T_1 == 8'hA2 & write_0_en];	// <stdin>:6285:13, :6286:13, :6287:13, :6289:13, :6292:9
      Register_inst163 <= _T_165[_T_1 == 8'hA3 & write_0_en];	// <stdin>:6300:13, :6301:13, :6302:13, :6304:13, :6307:9
      Register_inst164 <= _T_166[_T_1 == 8'hA4 & write_0_en];	// <stdin>:6315:13, :6316:13, :6317:13, :6319:13, :6322:9
      Register_inst165 <= _T_167[_T_1 == 8'hA5 & write_0_en];	// <stdin>:6330:13, :6331:13, :6332:13, :6334:13, :6337:9
      Register_inst166 <= _T_168[_T_1 == 8'hA6 & write_0_en];	// <stdin>:6345:13, :6346:13, :6347:13, :6349:13, :6352:9
      Register_inst167 <= _T_169[_T_1 == 8'hA7 & write_0_en];	// <stdin>:6360:13, :6361:13, :6362:13, :6364:13, :6367:9
      Register_inst168 <= _T_170[_T_1 == 8'hA8 & write_0_en];	// <stdin>:6375:13, :6376:13, :6377:13, :6379:13, :6382:9
      Register_inst169 <= _T_171[_T_1 == 8'hA9 & write_0_en];	// <stdin>:6390:13, :6391:13, :6392:13, :6394:13, :6397:9
      Register_inst170 <= _T_172[_T_1 == 8'hAA & write_0_en];	// <stdin>:6405:13, :6406:13, :6407:13, :6409:13, :6412:9
      Register_inst171 <= _T_173[_T_1 == 8'hAB & write_0_en];	// <stdin>:6420:13, :6421:13, :6422:13, :6424:13, :6427:9
      Register_inst172 <= _T_174[_T_1 == 8'hAC & write_0_en];	// <stdin>:6435:13, :6436:13, :6437:13, :6439:13, :6442:9
      Register_inst173 <= _T_175[_T_1 == 8'hAD & write_0_en];	// <stdin>:6450:13, :6451:13, :6452:13, :6454:13, :6457:9
      Register_inst174 <= _T_176[_T_1 == 8'hAE & write_0_en];	// <stdin>:6465:13, :6466:13, :6467:13, :6469:13, :6472:9
      Register_inst175 <= _T_177[_T_1 == 8'hAF & write_0_en];	// <stdin>:6480:13, :6481:13, :6482:13, :6484:13, :6487:9
      Register_inst176 <= _T_178[_T_1 == 8'hB0 & write_0_en];	// <stdin>:6495:13, :6496:13, :6497:13, :6499:13, :6502:9
      Register_inst177 <= _T_179[_T_1 == 8'hB1 & write_0_en];	// <stdin>:6510:13, :6511:13, :6512:13, :6514:13, :6517:9
      Register_inst178 <= _T_180[_T_1 == 8'hB2 & write_0_en];	// <stdin>:6525:13, :6526:13, :6527:13, :6529:13, :6532:9
      Register_inst179 <= _T_181[_T_1 == 8'hB3 & write_0_en];	// <stdin>:6540:13, :6541:13, :6542:13, :6544:13, :6547:9
      Register_inst180 <= _T_182[_T_1 == 8'hB4 & write_0_en];	// <stdin>:6555:13, :6556:13, :6557:13, :6559:13, :6562:9
      Register_inst181 <= _T_183[_T_1 == 8'hB5 & write_0_en];	// <stdin>:6570:13, :6571:13, :6572:13, :6574:13, :6577:9
      Register_inst182 <= _T_184[_T_1 == 8'hB6 & write_0_en];	// <stdin>:6585:13, :6586:13, :6587:13, :6589:13, :6592:9
      Register_inst183 <= _T_185[_T_1 == 8'hB7 & write_0_en];	// <stdin>:6600:13, :6601:13, :6602:13, :6604:13, :6607:9
      Register_inst184 <= _T_186[_T_1 == 8'hB8 & write_0_en];	// <stdin>:6615:13, :6616:13, :6617:13, :6619:13, :6622:9
      Register_inst185 <= _T_187[_T_1 == 8'hB9 & write_0_en];	// <stdin>:6630:13, :6631:13, :6632:13, :6634:13, :6637:9
      Register_inst186 <= _T_188[_T_1 == 8'hBA & write_0_en];	// <stdin>:6645:13, :6646:13, :6647:13, :6649:13, :6652:9
      Register_inst187 <= _T_189[_T_1 == 8'hBB & write_0_en];	// <stdin>:6660:13, :6661:13, :6662:13, :6664:13, :6667:9
      Register_inst188 <= _T_190[_T_1 == 8'hBC & write_0_en];	// <stdin>:6675:13, :6676:13, :6677:13, :6679:13, :6682:9
      Register_inst189 <= _T_191[_T_1 == 8'hBD & write_0_en];	// <stdin>:6690:13, :6691:13, :6692:13, :6694:13, :6697:9
      Register_inst190 <= _T_192[_T_1 == 8'hBE & write_0_en];	// <stdin>:6705:13, :6706:13, :6707:13, :6709:13, :6712:9
      Register_inst191 <= _T_193[_T_1 == 8'hBF & write_0_en];	// <stdin>:6720:13, :6721:13, :6722:13, :6724:13, :6727:9
      Register_inst192 <= _T_194[_T_1 == 8'hC0 & write_0_en];	// <stdin>:6735:13, :6736:13, :6737:13, :6739:13, :6742:9
      Register_inst193 <= _T_195[_T_1 == 8'hC1 & write_0_en];	// <stdin>:6750:13, :6751:13, :6752:13, :6754:13, :6757:9
      Register_inst194 <= _T_196[_T_1 == 8'hC2 & write_0_en];	// <stdin>:6765:13, :6766:13, :6767:13, :6769:13, :6772:9
      Register_inst195 <= _T_197[_T_1 == 8'hC3 & write_0_en];	// <stdin>:6780:13, :6781:13, :6782:13, :6784:13, :6787:9
      Register_inst196 <= _T_198[_T_1 == 8'hC4 & write_0_en];	// <stdin>:6795:13, :6796:13, :6797:13, :6799:13, :6802:9
      Register_inst197 <= _T_199[_T_1 == 8'hC5 & write_0_en];	// <stdin>:6810:13, :6811:13, :6812:13, :6814:13, :6817:9
      Register_inst198 <= _T_200[_T_1 == 8'hC6 & write_0_en];	// <stdin>:6825:13, :6826:13, :6827:13, :6829:13, :6832:9
      Register_inst199 <= _T_201[_T_1 == 8'hC7 & write_0_en];	// <stdin>:6840:13, :6841:13, :6842:13, :6844:13, :6847:9
      Register_inst200 <= _T_202[_T_1 == 8'hC8 & write_0_en];	// <stdin>:6855:13, :6856:13, :6857:13, :6859:13, :6862:9
      Register_inst201 <= _T_203[_T_1 == 8'hC9 & write_0_en];	// <stdin>:6870:13, :6871:13, :6872:13, :6874:13, :6877:9
      Register_inst202 <= _T_204[_T_1 == 8'hCA & write_0_en];	// <stdin>:6885:13, :6886:13, :6887:13, :6889:13, :6892:9
      Register_inst203 <= _T_205[_T_1 == 8'hCB & write_0_en];	// <stdin>:6900:13, :6901:13, :6902:13, :6904:13, :6907:9
      Register_inst204 <= _T_206[_T_1 == 8'hCC & write_0_en];	// <stdin>:6915:13, :6916:13, :6917:13, :6919:13, :6922:9
      Register_inst205 <= _T_207[_T_1 == 8'hCD & write_0_en];	// <stdin>:6930:13, :6931:13, :6932:13, :6934:13, :6937:9
      Register_inst206 <= _T_208[_T_1 == 8'hCE & write_0_en];	// <stdin>:6945:13, :6946:13, :6947:13, :6949:13, :6952:9
      Register_inst207 <= _T_209[_T_1 == 8'hCF & write_0_en];	// <stdin>:6960:13, :6961:13, :6962:13, :6964:13, :6967:9
      Register_inst208 <= _T_210[_T_1 == 8'hD0 & write_0_en];	// <stdin>:6975:13, :6976:13, :6977:13, :6979:13, :6982:9
      Register_inst209 <= _T_211[_T_1 == 8'hD1 & write_0_en];	// <stdin>:6990:13, :6991:13, :6992:13, :6994:13, :6997:9
      Register_inst210 <= _T_212[_T_1 == 8'hD2 & write_0_en];	// <stdin>:7005:13, :7006:13, :7007:13, :7009:13, :7012:9
      Register_inst211 <= _T_213[_T_1 == 8'hD3 & write_0_en];	// <stdin>:7020:13, :7021:13, :7022:13, :7024:13, :7027:9
      Register_inst212 <= _T_214[_T_1 == 8'hD4 & write_0_en];	// <stdin>:7035:13, :7036:13, :7037:13, :7039:13, :7042:9
      Register_inst213 <= _T_215[_T_1 == 8'hD5 & write_0_en];	// <stdin>:7050:13, :7051:13, :7052:13, :7054:13, :7057:9
      Register_inst214 <= _T_216[_T_1 == 8'hD6 & write_0_en];	// <stdin>:7065:13, :7066:13, :7067:13, :7069:13, :7072:9
      Register_inst215 <= _T_217[_T_1 == 8'hD7 & write_0_en];	// <stdin>:7080:13, :7081:13, :7082:13, :7084:13, :7087:9
      Register_inst216 <= _T_218[_T_1 == 8'hD8 & write_0_en];	// <stdin>:7095:13, :7096:13, :7097:13, :7099:13, :7102:9
      Register_inst217 <= _T_219[_T_1 == 8'hD9 & write_0_en];	// <stdin>:7110:13, :7111:13, :7112:13, :7114:13, :7117:9
      Register_inst218 <= _T_220[_T_1 == 8'hDA & write_0_en];	// <stdin>:7125:13, :7126:13, :7127:13, :7129:13, :7132:9
      Register_inst219 <= _T_221[_T_1 == 8'hDB & write_0_en];	// <stdin>:7140:13, :7141:13, :7142:13, :7144:13, :7147:9
      Register_inst220 <= _T_222[_T_1 == 8'hDC & write_0_en];	// <stdin>:7155:13, :7156:13, :7157:13, :7159:13, :7162:9
      Register_inst221 <= _T_223[_T_1 == 8'hDD & write_0_en];	// <stdin>:7170:13, :7171:13, :7172:13, :7174:13, :7177:9
      Register_inst222 <= _T_224[_T_1 == 8'hDE & write_0_en];	// <stdin>:7185:13, :7186:13, :7187:13, :7189:13, :7192:9
      Register_inst223 <= _T_225[_T_1 == 8'hDF & write_0_en];	// <stdin>:7200:13, :7201:13, :7202:13, :7204:13, :7207:9
      Register_inst224 <= _T_226[_T_1 == 8'hE0 & write_0_en];	// <stdin>:7215:13, :7216:13, :7217:13, :7219:13, :7222:9
      Register_inst225 <= _T_227[_T_1 == 8'hE1 & write_0_en];	// <stdin>:7230:13, :7231:13, :7232:13, :7234:13, :7237:9
      Register_inst226 <= _T_228[_T_1 == 8'hE2 & write_0_en];	// <stdin>:7245:13, :7246:13, :7247:13, :7249:13, :7252:9
      Register_inst227 <= _T_229[_T_1 == 8'hE3 & write_0_en];	// <stdin>:7260:13, :7261:13, :7262:13, :7264:13, :7267:9
      Register_inst228 <= _T_230[_T_1 == 8'hE4 & write_0_en];	// <stdin>:7275:13, :7276:13, :7277:13, :7279:13, :7282:9
      Register_inst229 <= _T_231[_T_1 == 8'hE5 & write_0_en];	// <stdin>:7290:13, :7291:13, :7292:13, :7294:13, :7297:9
      Register_inst230 <= _T_232[_T_1 == 8'hE6 & write_0_en];	// <stdin>:7305:13, :7306:13, :7307:13, :7309:13, :7312:9
      Register_inst231 <= _T_233[_T_1 == 8'hE7 & write_0_en];	// <stdin>:7320:13, :7321:13, :7322:13, :7324:13, :7327:9
      Register_inst232 <= _T_234[_T_1 == 8'hE8 & write_0_en];	// <stdin>:7335:13, :7336:13, :7337:13, :7339:13, :7342:9
      Register_inst233 <= _T_235[_T_1 == 8'hE9 & write_0_en];	// <stdin>:7350:13, :7351:13, :7352:13, :7354:13, :7357:9
      Register_inst234 <= _T_236[_T_1 == 8'hEA & write_0_en];	// <stdin>:7365:13, :7366:13, :7367:13, :7369:13, :7372:9
      Register_inst235 <= _T_237[_T_1 == 8'hEB & write_0_en];	// <stdin>:7380:13, :7381:13, :7382:13, :7384:13, :7387:9
      Register_inst236 <= _T_238[_T_1 == 8'hEC & write_0_en];	// <stdin>:7395:13, :7396:13, :7397:13, :7399:13, :7402:9
      Register_inst237 <= _T_239[_T_1 == 8'hED & write_0_en];	// <stdin>:7410:13, :7411:13, :7412:13, :7414:13, :7417:9
      Register_inst238 <= _T_240[_T_1 == 8'hEE & write_0_en];	// <stdin>:7425:13, :7426:13, :7427:13, :7429:13, :7432:9
      Register_inst239 <= _T_241[_T_1 == 8'hEF & write_0_en];	// <stdin>:7440:13, :7441:13, :7442:13, :7444:13, :7447:9
      Register_inst240 <= _T_242[_T_1 == 8'hF0 & write_0_en];	// <stdin>:7455:13, :7456:13, :7457:13, :7459:13, :7462:9
      Register_inst241 <= _T_243[_T_1 == 8'hF1 & write_0_en];	// <stdin>:7470:13, :7471:13, :7472:13, :7474:13, :7477:9
      Register_inst242 <= _T_244[_T_1 == 8'hF2 & write_0_en];	// <stdin>:7485:13, :7486:13, :7487:13, :7489:13, :7492:9
      Register_inst243 <= _T_245[_T_1 == 8'hF3 & write_0_en];	// <stdin>:7500:13, :7501:13, :7502:13, :7504:13, :7507:9
      Register_inst244 <= _T_246[_T_1 == 8'hF4 & write_0_en];	// <stdin>:7515:13, :7516:13, :7517:13, :7519:13, :7522:9
      Register_inst245 <= _T_247[_T_1 == 8'hF5 & write_0_en];	// <stdin>:7530:13, :7531:13, :7532:13, :7534:13, :7537:9
      Register_inst246 <= _T_248[_T_1 == 8'hF6 & write_0_en];	// <stdin>:7545:13, :7546:13, :7547:13, :7549:13, :7552:9
      Register_inst247 <= _T_249[_T_1 == 8'hF7 & write_0_en];	// <stdin>:7560:13, :7561:13, :7562:13, :7564:13, :7567:9
      Register_inst248 <= _T_250[_T_1 == 8'hF8 & write_0_en];	// <stdin>:7575:13, :7576:13, :7577:13, :7579:13, :7582:9
      Register_inst249 <= _T_251[_T_1 == 8'hF9 & write_0_en];	// <stdin>:7590:13, :7591:13, :7592:13, :7594:13, :7597:9
      Register_inst250 <= _T_252[_T_1 == 8'hFA & write_0_en];	// <stdin>:7605:13, :7606:13, :7607:13, :7609:13, :7612:9
      Register_inst251 <= _T_253[_T_1 == 8'hFB & write_0_en];	// <stdin>:7620:13, :7621:13, :7622:13, :7624:13, :7627:9
      Register_inst252 <= _T_254[_T_1 == 8'hFC & write_0_en];	// <stdin>:7635:13, :7636:13, :7637:13, :7639:13, :7642:9
      Register_inst253 <= _T_255[_T_1 == 8'hFD & write_0_en];	// <stdin>:7650:13, :7651:13, :7652:13, :7654:13, :7657:9
      Register_inst254 <= _T_256[_T_1 == 8'hFE & write_0_en];	// <stdin>:7665:13, :7666:13, :7667:13, :7669:13, :7672:9
      Register_inst255 <= _T_257[&_T_1 & write_0_en];	// <stdin>:7681:13, :7682:13, :7684:13, :7687:9
    end
  end // always_ff @(posedge or posedge)
  initial begin	// <stdin>:7691:5
    Register_inst0 = 32'h0;	// <stdin>:3865:10, :3867:9
    Register_inst1 = 32'h0;	// <stdin>:3865:10, :3882:9
    Register_inst2 = 32'h0;	// <stdin>:3865:10, :3897:9
    Register_inst3 = 32'h0;	// <stdin>:3865:10, :3912:9
    Register_inst4 = 32'h0;	// <stdin>:3865:10, :3927:9
    Register_inst5 = 32'h0;	// <stdin>:3865:10, :3942:9
    Register_inst6 = 32'h0;	// <stdin>:3865:10, :3957:9
    Register_inst7 = 32'h0;	// <stdin>:3865:10, :3972:9
    Register_inst8 = 32'h0;	// <stdin>:3865:10, :3987:9
    Register_inst9 = 32'h0;	// <stdin>:3865:10, :4002:9
    Register_inst10 = 32'h0;	// <stdin>:3865:10, :4017:9
    Register_inst11 = 32'h0;	// <stdin>:3865:10, :4032:9
    Register_inst12 = 32'h0;	// <stdin>:3865:10, :4047:9
    Register_inst13 = 32'h0;	// <stdin>:3865:10, :4062:9
    Register_inst14 = 32'h0;	// <stdin>:3865:10, :4077:9
    Register_inst15 = 32'h0;	// <stdin>:3865:10, :4092:9
    Register_inst16 = 32'h0;	// <stdin>:3865:10, :4107:9
    Register_inst17 = 32'h0;	// <stdin>:3865:10, :4122:9
    Register_inst18 = 32'h0;	// <stdin>:3865:10, :4137:9
    Register_inst19 = 32'h0;	// <stdin>:3865:10, :4152:9
    Register_inst20 = 32'h0;	// <stdin>:3865:10, :4167:9
    Register_inst21 = 32'h0;	// <stdin>:3865:10, :4182:9
    Register_inst22 = 32'h0;	// <stdin>:3865:10, :4197:9
    Register_inst23 = 32'h0;	// <stdin>:3865:10, :4212:9
    Register_inst24 = 32'h0;	// <stdin>:3865:10, :4227:9
    Register_inst25 = 32'h0;	// <stdin>:3865:10, :4242:9
    Register_inst26 = 32'h0;	// <stdin>:3865:10, :4257:9
    Register_inst27 = 32'h0;	// <stdin>:3865:10, :4272:9
    Register_inst28 = 32'h0;	// <stdin>:3865:10, :4287:9
    Register_inst29 = 32'h0;	// <stdin>:3865:10, :4302:9
    Register_inst30 = 32'h0;	// <stdin>:3865:10, :4317:9
    Register_inst31 = 32'h0;	// <stdin>:3865:10, :4332:9
    Register_inst32 = 32'h0;	// <stdin>:3865:10, :4347:9
    Register_inst33 = 32'h0;	// <stdin>:3865:10, :4362:9
    Register_inst34 = 32'h0;	// <stdin>:3865:10, :4377:9
    Register_inst35 = 32'h0;	// <stdin>:3865:10, :4392:9
    Register_inst36 = 32'h0;	// <stdin>:3865:10, :4407:9
    Register_inst37 = 32'h0;	// <stdin>:3865:10, :4422:9
    Register_inst38 = 32'h0;	// <stdin>:3865:10, :4437:9
    Register_inst39 = 32'h0;	// <stdin>:3865:10, :4452:9
    Register_inst40 = 32'h0;	// <stdin>:3865:10, :4467:9
    Register_inst41 = 32'h0;	// <stdin>:3865:10, :4482:9
    Register_inst42 = 32'h0;	// <stdin>:3865:10, :4497:9
    Register_inst43 = 32'h0;	// <stdin>:3865:10, :4512:9
    Register_inst44 = 32'h0;	// <stdin>:3865:10, :4527:9
    Register_inst45 = 32'h0;	// <stdin>:3865:10, :4542:9
    Register_inst46 = 32'h0;	// <stdin>:3865:10, :4557:9
    Register_inst47 = 32'h0;	// <stdin>:3865:10, :4572:9
    Register_inst48 = 32'h0;	// <stdin>:3865:10, :4587:9
    Register_inst49 = 32'h0;	// <stdin>:3865:10, :4602:9
    Register_inst50 = 32'h0;	// <stdin>:3865:10, :4617:9
    Register_inst51 = 32'h0;	// <stdin>:3865:10, :4632:9
    Register_inst52 = 32'h0;	// <stdin>:3865:10, :4647:9
    Register_inst53 = 32'h0;	// <stdin>:3865:10, :4662:9
    Register_inst54 = 32'h0;	// <stdin>:3865:10, :4677:9
    Register_inst55 = 32'h0;	// <stdin>:3865:10, :4692:9
    Register_inst56 = 32'h0;	// <stdin>:3865:10, :4707:9
    Register_inst57 = 32'h0;	// <stdin>:3865:10, :4722:9
    Register_inst58 = 32'h0;	// <stdin>:3865:10, :4737:9
    Register_inst59 = 32'h0;	// <stdin>:3865:10, :4752:9
    Register_inst60 = 32'h0;	// <stdin>:3865:10, :4767:9
    Register_inst61 = 32'h0;	// <stdin>:3865:10, :4782:9
    Register_inst62 = 32'h0;	// <stdin>:3865:10, :4797:9
    Register_inst63 = 32'h0;	// <stdin>:3865:10, :4812:9
    Register_inst64 = 32'h0;	// <stdin>:3865:10, :4827:9
    Register_inst65 = 32'h0;	// <stdin>:3865:10, :4842:9
    Register_inst66 = 32'h0;	// <stdin>:3865:10, :4857:9
    Register_inst67 = 32'h0;	// <stdin>:3865:10, :4872:9
    Register_inst68 = 32'h0;	// <stdin>:3865:10, :4887:9
    Register_inst69 = 32'h0;	// <stdin>:3865:10, :4902:9
    Register_inst70 = 32'h0;	// <stdin>:3865:10, :4917:9
    Register_inst71 = 32'h0;	// <stdin>:3865:10, :4932:9
    Register_inst72 = 32'h0;	// <stdin>:3865:10, :4947:9
    Register_inst73 = 32'h0;	// <stdin>:3865:10, :4962:9
    Register_inst74 = 32'h0;	// <stdin>:3865:10, :4977:9
    Register_inst75 = 32'h0;	// <stdin>:3865:10, :4992:9
    Register_inst76 = 32'h0;	// <stdin>:3865:10, :5007:9
    Register_inst77 = 32'h0;	// <stdin>:3865:10, :5022:9
    Register_inst78 = 32'h0;	// <stdin>:3865:10, :5037:9
    Register_inst79 = 32'h0;	// <stdin>:3865:10, :5052:9
    Register_inst80 = 32'h0;	// <stdin>:3865:10, :5067:9
    Register_inst81 = 32'h0;	// <stdin>:3865:10, :5082:9
    Register_inst82 = 32'h0;	// <stdin>:3865:10, :5097:9
    Register_inst83 = 32'h0;	// <stdin>:3865:10, :5112:9
    Register_inst84 = 32'h0;	// <stdin>:3865:10, :5127:9
    Register_inst85 = 32'h0;	// <stdin>:3865:10, :5142:9
    Register_inst86 = 32'h0;	// <stdin>:3865:10, :5157:9
    Register_inst87 = 32'h0;	// <stdin>:3865:10, :5172:9
    Register_inst88 = 32'h0;	// <stdin>:3865:10, :5187:9
    Register_inst89 = 32'h0;	// <stdin>:3865:10, :5202:9
    Register_inst90 = 32'h0;	// <stdin>:3865:10, :5217:9
    Register_inst91 = 32'h0;	// <stdin>:3865:10, :5232:9
    Register_inst92 = 32'h0;	// <stdin>:3865:10, :5247:9
    Register_inst93 = 32'h0;	// <stdin>:3865:10, :5262:9
    Register_inst94 = 32'h0;	// <stdin>:3865:10, :5277:9
    Register_inst95 = 32'h0;	// <stdin>:3865:10, :5292:9
    Register_inst96 = 32'h0;	// <stdin>:3865:10, :5307:9
    Register_inst97 = 32'h0;	// <stdin>:3865:10, :5322:9
    Register_inst98 = 32'h0;	// <stdin>:3865:10, :5337:9
    Register_inst99 = 32'h0;	// <stdin>:3865:10, :5352:9
    Register_inst100 = 32'h0;	// <stdin>:3865:10, :5367:9
    Register_inst101 = 32'h0;	// <stdin>:3865:10, :5382:9
    Register_inst102 = 32'h0;	// <stdin>:3865:10, :5397:9
    Register_inst103 = 32'h0;	// <stdin>:3865:10, :5412:9
    Register_inst104 = 32'h0;	// <stdin>:3865:10, :5427:9
    Register_inst105 = 32'h0;	// <stdin>:3865:10, :5442:9
    Register_inst106 = 32'h0;	// <stdin>:3865:10, :5457:9
    Register_inst107 = 32'h0;	// <stdin>:3865:10, :5472:9
    Register_inst108 = 32'h0;	// <stdin>:3865:10, :5487:9
    Register_inst109 = 32'h0;	// <stdin>:3865:10, :5502:9
    Register_inst110 = 32'h0;	// <stdin>:3865:10, :5517:9
    Register_inst111 = 32'h0;	// <stdin>:3865:10, :5532:9
    Register_inst112 = 32'h0;	// <stdin>:3865:10, :5547:9
    Register_inst113 = 32'h0;	// <stdin>:3865:10, :5562:9
    Register_inst114 = 32'h0;	// <stdin>:3865:10, :5577:9
    Register_inst115 = 32'h0;	// <stdin>:3865:10, :5592:9
    Register_inst116 = 32'h0;	// <stdin>:3865:10, :5607:9
    Register_inst117 = 32'h0;	// <stdin>:3865:10, :5622:9
    Register_inst118 = 32'h0;	// <stdin>:3865:10, :5637:9
    Register_inst119 = 32'h0;	// <stdin>:3865:10, :5652:9
    Register_inst120 = 32'h0;	// <stdin>:3865:10, :5667:9
    Register_inst121 = 32'h0;	// <stdin>:3865:10, :5682:9
    Register_inst122 = 32'h0;	// <stdin>:3865:10, :5697:9
    Register_inst123 = 32'h0;	// <stdin>:3865:10, :5712:9
    Register_inst124 = 32'h0;	// <stdin>:3865:10, :5727:9
    Register_inst125 = 32'h0;	// <stdin>:3865:10, :5742:9
    Register_inst126 = 32'h0;	// <stdin>:3865:10, :5757:9
    Register_inst127 = 32'h0;	// <stdin>:3865:10, :5772:9
    Register_inst128 = 32'h0;	// <stdin>:3865:10, :5787:9
    Register_inst129 = 32'h0;	// <stdin>:3865:10, :5802:9
    Register_inst130 = 32'h0;	// <stdin>:3865:10, :5817:9
    Register_inst131 = 32'h0;	// <stdin>:3865:10, :5832:9
    Register_inst132 = 32'h0;	// <stdin>:3865:10, :5847:9
    Register_inst133 = 32'h0;	// <stdin>:3865:10, :5862:9
    Register_inst134 = 32'h0;	// <stdin>:3865:10, :5877:9
    Register_inst135 = 32'h0;	// <stdin>:3865:10, :5892:9
    Register_inst136 = 32'h0;	// <stdin>:3865:10, :5907:9
    Register_inst137 = 32'h0;	// <stdin>:3865:10, :5922:9
    Register_inst138 = 32'h0;	// <stdin>:3865:10, :5937:9
    Register_inst139 = 32'h0;	// <stdin>:3865:10, :5952:9
    Register_inst140 = 32'h0;	// <stdin>:3865:10, :5967:9
    Register_inst141 = 32'h0;	// <stdin>:3865:10, :5982:9
    Register_inst142 = 32'h0;	// <stdin>:3865:10, :5997:9
    Register_inst143 = 32'h0;	// <stdin>:3865:10, :6012:9
    Register_inst144 = 32'h0;	// <stdin>:3865:10, :6027:9
    Register_inst145 = 32'h0;	// <stdin>:3865:10, :6042:9
    Register_inst146 = 32'h0;	// <stdin>:3865:10, :6057:9
    Register_inst147 = 32'h0;	// <stdin>:3865:10, :6072:9
    Register_inst148 = 32'h0;	// <stdin>:3865:10, :6087:9
    Register_inst149 = 32'h0;	// <stdin>:3865:10, :6102:9
    Register_inst150 = 32'h0;	// <stdin>:3865:10, :6117:9
    Register_inst151 = 32'h0;	// <stdin>:3865:10, :6132:9
    Register_inst152 = 32'h0;	// <stdin>:3865:10, :6147:9
    Register_inst153 = 32'h0;	// <stdin>:3865:10, :6162:9
    Register_inst154 = 32'h0;	// <stdin>:3865:10, :6177:9
    Register_inst155 = 32'h0;	// <stdin>:3865:10, :6192:9
    Register_inst156 = 32'h0;	// <stdin>:3865:10, :6207:9
    Register_inst157 = 32'h0;	// <stdin>:3865:10, :6222:9
    Register_inst158 = 32'h0;	// <stdin>:3865:10, :6237:9
    Register_inst159 = 32'h0;	// <stdin>:3865:10, :6252:9
    Register_inst160 = 32'h0;	// <stdin>:3865:10, :6267:9
    Register_inst161 = 32'h0;	// <stdin>:3865:10, :6282:9
    Register_inst162 = 32'h0;	// <stdin>:3865:10, :6297:9
    Register_inst163 = 32'h0;	// <stdin>:3865:10, :6312:9
    Register_inst164 = 32'h0;	// <stdin>:3865:10, :6327:9
    Register_inst165 = 32'h0;	// <stdin>:3865:10, :6342:9
    Register_inst166 = 32'h0;	// <stdin>:3865:10, :6357:9
    Register_inst167 = 32'h0;	// <stdin>:3865:10, :6372:9
    Register_inst168 = 32'h0;	// <stdin>:3865:10, :6387:9
    Register_inst169 = 32'h0;	// <stdin>:3865:10, :6402:9
    Register_inst170 = 32'h0;	// <stdin>:3865:10, :6417:9
    Register_inst171 = 32'h0;	// <stdin>:3865:10, :6432:9
    Register_inst172 = 32'h0;	// <stdin>:3865:10, :6447:9
    Register_inst173 = 32'h0;	// <stdin>:3865:10, :6462:9
    Register_inst174 = 32'h0;	// <stdin>:3865:10, :6477:9
    Register_inst175 = 32'h0;	// <stdin>:3865:10, :6492:9
    Register_inst176 = 32'h0;	// <stdin>:3865:10, :6507:9
    Register_inst177 = 32'h0;	// <stdin>:3865:10, :6522:9
    Register_inst178 = 32'h0;	// <stdin>:3865:10, :6537:9
    Register_inst179 = 32'h0;	// <stdin>:3865:10, :6552:9
    Register_inst180 = 32'h0;	// <stdin>:3865:10, :6567:9
    Register_inst181 = 32'h0;	// <stdin>:3865:10, :6582:9
    Register_inst182 = 32'h0;	// <stdin>:3865:10, :6597:9
    Register_inst183 = 32'h0;	// <stdin>:3865:10, :6612:9
    Register_inst184 = 32'h0;	// <stdin>:3865:10, :6627:9
    Register_inst185 = 32'h0;	// <stdin>:3865:10, :6642:9
    Register_inst186 = 32'h0;	// <stdin>:3865:10, :6657:9
    Register_inst187 = 32'h0;	// <stdin>:3865:10, :6672:9
    Register_inst188 = 32'h0;	// <stdin>:3865:10, :6687:9
    Register_inst189 = 32'h0;	// <stdin>:3865:10, :6702:9
    Register_inst190 = 32'h0;	// <stdin>:3865:10, :6717:9
    Register_inst191 = 32'h0;	// <stdin>:3865:10, :6732:9
    Register_inst192 = 32'h0;	// <stdin>:3865:10, :6747:9
    Register_inst193 = 32'h0;	// <stdin>:3865:10, :6762:9
    Register_inst194 = 32'h0;	// <stdin>:3865:10, :6777:9
    Register_inst195 = 32'h0;	// <stdin>:3865:10, :6792:9
    Register_inst196 = 32'h0;	// <stdin>:3865:10, :6807:9
    Register_inst197 = 32'h0;	// <stdin>:3865:10, :6822:9
    Register_inst198 = 32'h0;	// <stdin>:3865:10, :6837:9
    Register_inst199 = 32'h0;	// <stdin>:3865:10, :6852:9
    Register_inst200 = 32'h0;	// <stdin>:3865:10, :6867:9
    Register_inst201 = 32'h0;	// <stdin>:3865:10, :6882:9
    Register_inst202 = 32'h0;	// <stdin>:3865:10, :6897:9
    Register_inst203 = 32'h0;	// <stdin>:3865:10, :6912:9
    Register_inst204 = 32'h0;	// <stdin>:3865:10, :6927:9
    Register_inst205 = 32'h0;	// <stdin>:3865:10, :6942:9
    Register_inst206 = 32'h0;	// <stdin>:3865:10, :6957:9
    Register_inst207 = 32'h0;	// <stdin>:3865:10, :6972:9
    Register_inst208 = 32'h0;	// <stdin>:3865:10, :6987:9
    Register_inst209 = 32'h0;	// <stdin>:3865:10, :7002:9
    Register_inst210 = 32'h0;	// <stdin>:3865:10, :7017:9
    Register_inst211 = 32'h0;	// <stdin>:3865:10, :7032:9
    Register_inst212 = 32'h0;	// <stdin>:3865:10, :7047:9
    Register_inst213 = 32'h0;	// <stdin>:3865:10, :7062:9
    Register_inst214 = 32'h0;	// <stdin>:3865:10, :7077:9
    Register_inst215 = 32'h0;	// <stdin>:3865:10, :7092:9
    Register_inst216 = 32'h0;	// <stdin>:3865:10, :7107:9
    Register_inst217 = 32'h0;	// <stdin>:3865:10, :7122:9
    Register_inst218 = 32'h0;	// <stdin>:3865:10, :7137:9
    Register_inst219 = 32'h0;	// <stdin>:3865:10, :7152:9
    Register_inst220 = 32'h0;	// <stdin>:3865:10, :7167:9
    Register_inst221 = 32'h0;	// <stdin>:3865:10, :7182:9
    Register_inst222 = 32'h0;	// <stdin>:3865:10, :7197:9
    Register_inst223 = 32'h0;	// <stdin>:3865:10, :7212:9
    Register_inst224 = 32'h0;	// <stdin>:3865:10, :7227:9
    Register_inst225 = 32'h0;	// <stdin>:3865:10, :7242:9
    Register_inst226 = 32'h0;	// <stdin>:3865:10, :7257:9
    Register_inst227 = 32'h0;	// <stdin>:3865:10, :7272:9
    Register_inst228 = 32'h0;	// <stdin>:3865:10, :7287:9
    Register_inst229 = 32'h0;	// <stdin>:3865:10, :7302:9
    Register_inst230 = 32'h0;	// <stdin>:3865:10, :7317:9
    Register_inst231 = 32'h0;	// <stdin>:3865:10, :7332:9
    Register_inst232 = 32'h0;	// <stdin>:3865:10, :7347:9
    Register_inst233 = 32'h0;	// <stdin>:3865:10, :7362:9
    Register_inst234 = 32'h0;	// <stdin>:3865:10, :7377:9
    Register_inst235 = 32'h0;	// <stdin>:3865:10, :7392:9
    Register_inst236 = 32'h0;	// <stdin>:3865:10, :7407:9
    Register_inst237 = 32'h0;	// <stdin>:3865:10, :7422:9
    Register_inst238 = 32'h0;	// <stdin>:3865:10, :7437:9
    Register_inst239 = 32'h0;	// <stdin>:3865:10, :7452:9
    Register_inst240 = 32'h0;	// <stdin>:3865:10, :7467:9
    Register_inst241 = 32'h0;	// <stdin>:3865:10, :7482:9
    Register_inst242 = 32'h0;	// <stdin>:3865:10, :7497:9
    Register_inst243 = 32'h0;	// <stdin>:3865:10, :7512:9
    Register_inst244 = 32'h0;	// <stdin>:3865:10, :7527:9
    Register_inst245 = 32'h0;	// <stdin>:3865:10, :7542:9
    Register_inst246 = 32'h0;	// <stdin>:3865:10, :7557:9
    Register_inst247 = 32'h0;	// <stdin>:3865:10, :7572:9
    Register_inst248 = 32'h0;	// <stdin>:3865:10, :7587:9
    Register_inst249 = 32'h0;	// <stdin>:3865:10, :7602:9
    Register_inst250 = 32'h0;	// <stdin>:3865:10, :7617:9
    Register_inst251 = 32'h0;	// <stdin>:3865:10, :7632:9
    Register_inst252 = 32'h0;	// <stdin>:3865:10, :7647:9
    Register_inst253 = 32'h0;	// <stdin>:3865:10, :7662:9
    Register_inst254 = 32'h0;	// <stdin>:3865:10, :7677:9
    Register_inst255 = 32'h0;	// <stdin>:3865:10, :7692:9
  end // initial
  wire [255:0][31:0] _T = {{Register_inst0}, {Register_inst1}, {Register_inst2}, {Register_inst3}, {Register_inst4},
                {Register_inst5}, {Register_inst6}, {Register_inst7}, {Register_inst8}, {Register_inst9},
                {Register_inst10}, {Register_inst11}, {Register_inst12}, {Register_inst13},
                {Register_inst14}, {Register_inst15}, {Register_inst16}, {Register_inst17},
                {Register_inst18}, {Register_inst19}, {Register_inst20}, {Register_inst21},
                {Register_inst22}, {Register_inst23}, {Register_inst24}, {Register_inst25},
                {Register_inst26}, {Register_inst27}, {Register_inst28}, {Register_inst29},
                {Register_inst30}, {Register_inst31}, {Register_inst32}, {Register_inst33},
                {Register_inst34}, {Register_inst35}, {Register_inst36}, {Register_inst37},
                {Register_inst38}, {Register_inst39}, {Register_inst40}, {Register_inst41},
                {Register_inst42}, {Register_inst43}, {Register_inst44}, {Register_inst45},
                {Register_inst46}, {Register_inst47}, {Register_inst48}, {Register_inst49},
                {Register_inst50}, {Register_inst51}, {Register_inst52}, {Register_inst53},
                {Register_inst54}, {Register_inst55}, {Register_inst56}, {Register_inst57},
                {Register_inst58}, {Register_inst59}, {Register_inst60}, {Register_inst61},
                {Register_inst62}, {Register_inst63}, {Register_inst64}, {Register_inst65},
                {Register_inst66}, {Register_inst67}, {Register_inst68}, {Register_inst69},
                {Register_inst70}, {Register_inst71}, {Register_inst72}, {Register_inst73},
                {Register_inst74}, {Register_inst75}, {Register_inst76}, {Register_inst77},
                {Register_inst78}, {Register_inst79}, {Register_inst80}, {Register_inst81},
                {Register_inst82}, {Register_inst83}, {Register_inst84}, {Register_inst85},
                {Register_inst86}, {Register_inst87}, {Register_inst88}, {Register_inst89},
                {Register_inst90}, {Register_inst91}, {Register_inst92}, {Register_inst93},
                {Register_inst94}, {Register_inst95}, {Register_inst96}, {Register_inst97},
                {Register_inst98}, {Register_inst99}, {Register_inst100}, {Register_inst101},
                {Register_inst102}, {Register_inst103}, {Register_inst104}, {Register_inst105},
                {Register_inst106}, {Register_inst107}, {Register_inst108}, {Register_inst109},
                {Register_inst110}, {Register_inst111}, {Register_inst112}, {Register_inst113},
                {Register_inst114}, {Register_inst115}, {Register_inst116}, {Register_inst117},
                {Register_inst118}, {Register_inst119}, {Register_inst120}, {Register_inst121},
                {Register_inst122}, {Register_inst123}, {Register_inst124}, {Register_inst125},
                {Register_inst126}, {Register_inst127}, {Register_inst128}, {Register_inst129},
                {Register_inst130}, {Register_inst131}, {Register_inst132}, {Register_inst133},
                {Register_inst134}, {Register_inst135}, {Register_inst136}, {Register_inst137},
                {Register_inst138}, {Register_inst139}, {Register_inst140}, {Register_inst141},
                {Register_inst142}, {Register_inst143}, {Register_inst144}, {Register_inst145},
                {Register_inst146}, {Register_inst147}, {Register_inst148}, {Register_inst149},
                {Register_inst150}, {Register_inst151}, {Register_inst152}, {Register_inst153},
                {Register_inst154}, {Register_inst155}, {Register_inst156}, {Register_inst157},
                {Register_inst158}, {Register_inst159}, {Register_inst160}, {Register_inst161},
                {Register_inst162}, {Register_inst163}, {Register_inst164}, {Register_inst165},
                {Register_inst166}, {Register_inst167}, {Register_inst168}, {Register_inst169},
                {Register_inst170}, {Register_inst171}, {Register_inst172}, {Register_inst173},
                {Register_inst174}, {Register_inst175}, {Register_inst176}, {Register_inst177},
                {Register_inst178}, {Register_inst179}, {Register_inst180}, {Register_inst181},
                {Register_inst182}, {Register_inst183}, {Register_inst184}, {Register_inst185},
                {Register_inst186}, {Register_inst187}, {Register_inst188}, {Register_inst189},
                {Register_inst190}, {Register_inst191}, {Register_inst192}, {Register_inst193},
                {Register_inst194}, {Register_inst195}, {Register_inst196}, {Register_inst197},
                {Register_inst198}, {Register_inst199}, {Register_inst200}, {Register_inst201},
                {Register_inst202}, {Register_inst203}, {Register_inst204}, {Register_inst205},
                {Register_inst206}, {Register_inst207}, {Register_inst208}, {Register_inst209},
                {Register_inst210}, {Register_inst211}, {Register_inst212}, {Register_inst213},
                {Register_inst214}, {Register_inst215}, {Register_inst216}, {Register_inst217},
                {Register_inst218}, {Register_inst219}, {Register_inst220}, {Register_inst221},
                {Register_inst222}, {Register_inst223}, {Register_inst224}, {Register_inst225},
                {Register_inst226}, {Register_inst227}, {Register_inst228}, {Register_inst229},
                {Register_inst230}, {Register_inst231}, {Register_inst232}, {Register_inst233},
                {Register_inst234}, {Register_inst235}, {Register_inst236}, {Register_inst237},
                {Register_inst238}, {Register_inst239}, {Register_inst240}, {Register_inst241},
                {Register_inst242}, {Register_inst243}, {Register_inst244}, {Register_inst245},
                {Register_inst246}, {Register_inst247}, {Register_inst248}, {Register_inst249},
                {Register_inst250}, {Register_inst251}, {Register_inst252}, {Register_inst253},
                {Register_inst254}, {Register_inst255}};	// <stdin>:3869:10, :3884:11, :3899:11, :3914:11, :3929:11, :3944:11, :3959:11, :3974:11, :3989:11, :4004:11, :4019:11, :4034:11, :4049:11, :4064:11, :4079:12, :4094:12, :4109:12, :4124:12, :4139:12, :4154:12, :4169:12, :4184:12, :4199:12, :4214:12, :4229:12, :4244:12, :4259:12, :4274:12, :4289:12, :4304:12, :4319:12, :4334:12, :4349:12, :4364:12, :4379:12, :4394:12, :4409:12, :4424:12, :4439:12, :4454:12, :4469:12, :4484:12, :4499:12, :4514:12, :4529:12, :4544:12, :4559:12, :4574:12, :4589:12, :4604:12, :4619:12, :4634:12, :4649:12, :4664:12, :4679:12, :4694:12, :4709:12, :4724:12, :4739:12, :4754:12, :4769:12, :4784:12, :4799:12, :4814:12, :4829:12, :4844:12, :4859:12, :4874:12, :4889:12, :4904:12, :4919:12, :4934:12, :4949:12, :4964:12, :4979:12, :4994:12, :5009:12, :5024:12, :5039:12, :5054:12, :5069:12, :5084:12, :5099:12, :5114:12, :5129:12, :5144:12, :5159:12, :5174:12, :5189:12, :5204:12, :5219:12, :5234:12, :5249:12, :5264:12, :5279:12, :5294:12, :5309:12, :5324:12, :5339:12, :5354:12, :5369:12, :5384:12, :5399:12, :5414:12, :5429:12, :5444:12, :5459:12, :5474:12, :5489:12, :5504:12, :5519:12, :5534:12, :5549:12, :5564:12, :5579:12, :5594:12, :5609:12, :5624:12, :5639:12, :5654:12, :5669:12, :5684:12, :5699:12, :5714:12, :5729:12, :5744:12, :5759:12, :5774:12, :5789:12, :5804:12, :5819:12, :5834:12, :5849:12, :5864:12, :5879:12, :5894:12, :5909:12, :5924:12, :5939:12, :5954:12, :5969:12, :5984:12, :5999:13, :6014:13, :6029:13, :6044:13, :6059:13, :6074:13, :6089:13, :6104:13, :6119:13, :6134:13, :6149:13, :6164:13, :6179:13, :6194:13, :6209:13, :6224:13, :6239:13, :6254:13, :6269:13, :6284:13, :6299:13, :6314:13, :6329:13, :6344:13, :6359:13, :6374:13, :6389:13, :6404:13, :6419:13, :6434:13, :6449:13, :6464:13, :6479:13, :6494:13, :6509:13, :6524:13, :6539:13, :6554:13, :6569:13, :6584:13, :6599:13, :6614:13, :6629:13, :6644:13, :6659:13, :6674:13, :6689:13, :6704:13, :6719:13, :6734:13, :6749:13, :6764:13, :6779:13, :6794:13, :6809:13, :6824:13, :6839:13, :6854:13, :6869:13, :6884:13, :6899:13, :6914:13, :6929:13, :6944:13, :6959:13, :6974:13, :6989:13, :7004:13, :7019:13, :7034:13, :7049:13, :7064:13, :7079:13, :7094:13, :7109:13, :7124:13, :7139:13, :7154:13, :7169:13, :7184:13, :7199:13, :7214:13, :7229:13, :7244:13, :7259:13, :7274:13, :7289:13, :7304:13, :7319:13, :7334:13, :7349:13, :7364:13, :7379:13, :7394:13, :7409:13, :7424:13, :7439:13, :7454:13, :7469:13, :7484:13, :7499:13, :7514:13, :7529:13, :7544:13, :7559:13, :7574:13, :7589:13, :7604:13, :7619:13, :7634:13, :7649:13, :7664:13, :7679:13, :7694:13, :7695:13
  assign code_read_0_data = _T[code_read_0_addr];	// <stdin>:7696:13, :7697:5
endmodule

module Risc(	// <stdin>:7699:1
  input         is_write,
  input  [7:0]  write_addr,
  input  [31:0] write_data,
  input         boot, CLK, ASYNCRESET,
  output        valid,
  output [31:0] out);

  wire [31:0] _T;	// <stdin>:7840:12
  wire [31:0] file_file_read_0_data;	// <stdin>:7816:18
  wire [31:0] file_file_read_1_data;	// <stdin>:7816:18
  wire [31:0] code_code_read_0_data;	// <stdin>:7719:11
  reg  [7:0]  Register_inst0;	// <stdin>:7709:11

  always_ff @(posedge CLK) begin	// <stdin>:7710:5
    automatic logic [1:0][7:0] _T_11 = {{Register_inst0 + 8'h1}, {8'h0}};	// <stdin>:7702:10, :7703:10, :7704:10, :7705:10, :7717:10
    automatic logic [1:0][7:0] _T_12 = {{_T_11[boot]}, {Register_inst0}};	// <stdin>:7706:10, :7707:10, :7717:10

    Register_inst0 <= _T_12[is_write];	// <stdin>:7708:10, :7711:9
  end // always_ff @(posedge)
  initial	// <stdin>:7714:5
    Register_inst0 = 8'h0;	// <stdin>:7704:10, :7715:9
  wire struct packed {logic [31:0] data; logic [7:0] addr; } _T_0 = '{data: write_data, addr: write_addr};	// <stdin>:7718:11
  wire [1:0] _T_1 = {{1'h0}, {1'h1}};	// <stdin>:7700:10, :7701:10, :7731:11
  wire [1:0] _T_2 = {{_T_1[&(code_code_read_0_data[23:16])]}, {1'h0}};	// <stdin>:7700:10, :7719:11, :7728:11, :7730:11, :7732:11, :7734:11
  wire [1:0] _T_3 = {{_T_2[boot]}, {1'h0}};	// <stdin>:7700:10, :7735:11, :7737:11
  wire [1:0][31:0] _T_4 = {{32'h0}, {{24'h0, code_code_read_0_data[7:0]}}};	// <stdin>:7719:11, :7739:11, :7793:11, :7805:12
  wire struct packed {logic [31:0] data; logic [7:0] addr; } _T_5 = '{data: _T, addr: (code_code_read_0_data[23:16])};	// <stdin>:7719:11, :7809:12, :7810:12, :7840:12
  wire [1:0][31:0] _T_6 = {{file_file_read_0_data}, {32'h0}};	// <stdin>:7739:11, :7816:18, :7821:12
  wire [1:0][31:0] _T_7 = {{file_file_read_1_data}, {32'h0}};	// <stdin>:7739:11, :7816:18, :7827:12
  wire [1:0][31:0] _T_8 = {{_T_4[code_code_read_0_data[31:24] == 8'h1]}, {_T_6[code_code_read_0_data[15:8] == 8'h0] +
                _T_7[code_code_read_0_data[7:0] == 8'h0]}};	// <stdin>:7702:10, :7704:10, :7719:11, :7802:11, :7804:11, :7806:11, :7818:12, :7820:12, :7822:12, :7824:12, :7826:12, :7828:12, :7829:12, :7833:12
  wire [1:0][31:0] _T_9 = {{_T_8[code_code_read_0_data[31:24] == 8'h0]}, {32'h0}};	// <stdin>:7704:10, :7719:11, :7739:11, :7830:12, :7832:12, :7834:12, :7836:12
  wire [1:0][31:0] _T_10 = {{_T_9[boot]}, {32'h0}};	// <stdin>:7739:11, :7837:12, :7839:12
  assign _T = _T_10[is_write];	// <stdin>:7840:12
  code code (	// <stdin>:7719:11
    .CLK              (CLK),
    .ASYNCRESET       (ASYNCRESET),
    .code_read_0_addr (Register_inst0),	// <stdin>:7717:10
    .write_0          (_T_0),
    .write_0_en       (is_write),
    .code_read_0_data (code_code_read_0_data)
  );
  file file (	// <stdin>:7816:18
    .CLK              (CLK),
    .ASYNCRESET       (ASYNCRESET),
    .file_read_0_addr (code_code_read_0_data[15:8]),	// <stdin>:7719:11, :7807:12
    .file_read_1_addr (code_code_read_0_data[7:0]),	// <stdin>:7719:11, :7808:12
    .write_0          (_T_5),
    .write_0_en       (code_code_read_0_data[23:16] != 8'hFF),	// <stdin>:7719:11, :7729:11, :7811:12, :7813:12
    .file_read_0_data (file_file_read_0_data),
    .file_read_1_data (file_file_read_1_data)
  );
  assign valid = _T_3[is_write];	// <stdin>:7738:11, :7841:5
  assign out = _T;	// <stdin>:7840:12, :7841:5
endmodule

