module mod4 #(parameter KRATOS_INSTANCE_ID = 13'o7)
(
    input I
);

endmodule   // mod
