module return_py_tuple (input [1:0] I_0, output  O0, output  O1);
assign O0 = I_0[0];
assign O1 = I_0[1];
endmodule

