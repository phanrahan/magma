module mantle_slicesArrT__slices4220__t_0BitIn_1BitIn24 (
    input in_0__0,
    input [1:0] in_0__1,
    input in_1__0,
    input [1:0] in_1__1,
    input in_2__0,
    input [1:0] in_2__1,
    input in_3__0,
    input [1:0] in_3__1,
    output out0_0__0,
    output [1:0] out0_0__1,
    output out0_1__0,
    output [1:0] out0_1__1,
    output out1_0__0,
    output [1:0] out1_0__1,
    output out1_1__0,
    output [1:0] out1_1__1
);
assign out0_0__0 = in_2__0;
assign out0_0__1 = in_2__1;
assign out0_1__0 = in_3__0;
assign out0_1__1 = in_3__1;
assign out1_0__0 = in_0__0;
assign out1_0__1 = in_0__1;
assign out1_1__0 = in_1__0;
assign out1_1__1 = in_1__1;
endmodule

module mantle_liftArrT__t_0Bit_1Bit21 (
    input in__0,
    input [1:0] in__1,
    output out_0__0,
    output [1:0] out_0__1
);
assign out_0__0 = in__0;
assign out_0__1 = in__1;
endmodule

module mantle_concatNArrT__Ns22__t_child_0BitIn_1BitIn2 (
    input in0_0__0,
    input [1:0] in0_0__1,
    input in0_1__0,
    input [1:0] in0_1__1,
    input in1_0__0,
    input [1:0] in1_0__1,
    input in1_1__0,
    input [1:0] in1_1__1,
    output out_0__0,
    output [1:0] out_0__1,
    output out_1__0,
    output [1:0] out_1__1,
    output out_2__0,
    output [1:0] out_2__1,
    output out_3__0,
    output [1:0] out_3__1
);
assign out_0__0 = in0_0__0;
assign out_0__1 = in0_0__1;
assign out_1__0 = in0_1__0;
assign out_1__1 = in0_1__1;
assign out_2__0 = in1_0__0;
assign out_2__1 = in1_0__1;
assign out_3__0 = in1_1__0;
assign out_3__1 = in1_1__1;
endmodule

module mantle_concatNArrT__Ns1__t_child_0BitIn_1BitIn2 (
    input in0_0__0,
    input [1:0] in0_0__1,
    output out_0__0,
    output [1:0] out_0__1
);
assign out_0__0 = in0_0__0;
assign out_0__1 = in0_0__1;
endmodule

module mantle_concatNArrT__Ns13__t_child_0BitIn_1BitIn2 (
    input in0_0__0,
    input [1:0] in0_0__1,
    input in1_0__0,
    input [1:0] in1_0__1,
    input in1_1__0,
    input [1:0] in1_1__1,
    input in1_2__0,
    input [1:0] in1_2__1,
    output out_0__0,
    output [1:0] out_0__1,
    output out_1__0,
    output [1:0] out_1__1,
    output out_2__0,
    output [1:0] out_2__1,
    output out_3__0,
    output [1:0] out_3__1
);
assign out_0__0 = in0_0__0;
assign out_0__1 = in0_0__1;
assign out_1__0 = in1_0__0;
assign out_1__1 = in1_0__1;
assign out_2__0 = in1_1__0;
assign out_2__1 = in1_1__1;
assign out_3__0 = in1_2__0;
assign out_3__1 = in1_2__1;
endmodule

module mantle_concatNArrT__Ns12__t_child_0BitIn_1BitIn2 (
    input in0_0__0,
    input [1:0] in0_0__1,
    input in1_0__0,
    input [1:0] in1_0__1,
    input in1_1__0,
    input [1:0] in1_1__1,
    output out_0__0,
    output [1:0] out_0__1,
    output out_1__0,
    output [1:0] out_1__1,
    output out_2__0,
    output [1:0] out_2__1
);
assign out_0__0 = in0_0__0;
assign out_0__1 = in0_0__1;
assign out_1__0 = in1_0__0;
assign out_1__1 = in1_0__1;
assign out_2__0 = in1_1__0;
assign out_2__1 = in1_1__1;
endmodule

module mantle_concatNArrT__Ns11__t_child_0BitIn_1BitIn2 (
    input in0_0__0,
    input [1:0] in0_0__1,
    input in1_0__0,
    input [1:0] in1_0__1,
    output out_0__0,
    output [1:0] out_0__1,
    output out_1__0,
    output [1:0] out_1__1
);
assign out_0__0 = in0_0__0;
assign out_0__1 = in0_0__1;
assign out_1__0 = in1_0__0;
assign out_1__1 = in1_0__1;
endmodule

module Foo (
    input I_0__0,
    input [1:0] I_0__1,
    input I_1__0,
    input [1:0] I_1__1,
    input I_2__0,
    input [1:0] I_2__1,
    input I_3__0,
    input [1:0] I_3__1,
    output O0_0__0,
    output [1:0] O0_0__1,
    output O0_1__0,
    output [1:0] O0_1__1,
    output O0_2__0,
    output [1:0] O0_2__1,
    output O0_3__0,
    output [1:0] O0_3__1,
    output O1_0__0,
    output [1:0] O1_0__1,
    output O1_1__0,
    output [1:0] O1_1__1,
    output O1_2__0,
    output [1:0] O1_2__1,
    output O1_3__0,
    output [1:0] O1_3__1,
    output O2_0__0,
    output [1:0] O2_0__1,
    output O2_1__0,
    output [1:0] O2_1__1,
    output O2_2__0,
    output [1:0] O2_2__1,
    output O2_3__0,
    output [1:0] O2_3__1,
    output O3_0__0,
    output [1:0] O3_0__1,
    output O3_1__0,
    output [1:0] O3_1__1,
    output O3_2__0,
    output [1:0] O3_2__1,
    output O3_3__0,
    output [1:0] O3_3__1
);
wire ConcatN_inst0_out_0__0;
wire [1:0] ConcatN_inst0_out_0__1;
wire ConcatN_inst0_out_1__0;
wire [1:0] ConcatN_inst0_out_1__1;
wire ConcatN_inst0_out_2__0;
wire [1:0] ConcatN_inst0_out_2__1;
wire ConcatN_inst0_out_3__0;
wire [1:0] ConcatN_inst0_out_3__1;
wire ConcatN_inst1_out_0__0;
wire [1:0] ConcatN_inst1_out_0__1;
wire ConcatN_inst1_out_1__0;
wire [1:0] ConcatN_inst1_out_1__1;
wire ConcatN_inst1_out_2__0;
wire [1:0] ConcatN_inst1_out_2__1;
wire ConcatN_inst1_out_3__0;
wire [1:0] ConcatN_inst1_out_3__1;
wire ConcatN_inst2_out_0__0;
wire [1:0] ConcatN_inst2_out_0__1;
wire ConcatN_inst2_out_1__0;
wire [1:0] ConcatN_inst2_out_1__1;
wire ConcatN_inst2_out_2__0;
wire [1:0] ConcatN_inst2_out_2__1;
wire ConcatN_inst3_out_0__0;
wire [1:0] ConcatN_inst3_out_0__1;
wire ConcatN_inst3_out_1__0;
wire [1:0] ConcatN_inst3_out_1__1;
wire ConcatN_inst4_out_0__0;
wire [1:0] ConcatN_inst4_out_0__1;
wire ConcatN_inst5_out_0__0;
wire [1:0] ConcatN_inst5_out_0__1;
wire ConcatN_inst5_out_1__0;
wire [1:0] ConcatN_inst5_out_1__1;
wire ConcatN_inst5_out_2__0;
wire [1:0] ConcatN_inst5_out_2__1;
wire ConcatN_inst5_out_3__0;
wire [1:0] ConcatN_inst5_out_3__1;
wire Lift_inst0_out_0__0;
wire [1:0] Lift_inst0_out_0__1;
wire Lift_inst1_out_0__0;
wire [1:0] Lift_inst1_out_0__1;
wire Lift_inst2_out_0__0;
wire [1:0] Lift_inst2_out_0__1;
wire Lift_inst3_out_0__0;
wire [1:0] Lift_inst3_out_0__1;
wire SlicesBuilder_out0_0__0;
wire [1:0] SlicesBuilder_out0_0__1;
wire SlicesBuilder_out0_1__0;
wire [1:0] SlicesBuilder_out0_1__1;
wire SlicesBuilder_out1_0__0;
wire [1:0] SlicesBuilder_out1_0__1;
wire SlicesBuilder_out1_1__0;
wire [1:0] SlicesBuilder_out1_1__1;
mantle_concatNArrT__Ns22__t_child_0BitIn_1BitIn2 ConcatN_inst0 (
    .in0_0__0(SlicesBuilder_out0_0__0),
    .in0_0__1(SlicesBuilder_out0_0__1),
    .in0_1__0(SlicesBuilder_out0_1__0),
    .in0_1__1(SlicesBuilder_out0_1__1),
    .in1_0__0(SlicesBuilder_out1_0__0),
    .in1_0__1(SlicesBuilder_out1_0__1),
    .in1_1__0(SlicesBuilder_out1_1__0),
    .in1_1__1(SlicesBuilder_out1_1__1),
    .out_0__0(ConcatN_inst0_out_0__0),
    .out_0__1(ConcatN_inst0_out_0__1),
    .out_1__0(ConcatN_inst0_out_1__0),
    .out_1__1(ConcatN_inst0_out_1__1),
    .out_2__0(ConcatN_inst0_out_2__0),
    .out_2__1(ConcatN_inst0_out_2__1),
    .out_3__0(ConcatN_inst0_out_3__0),
    .out_3__1(ConcatN_inst0_out_3__1)
);
mantle_concatNArrT__Ns13__t_child_0BitIn_1BitIn2 ConcatN_inst1 (
    .in0_0__0(Lift_inst0_out_0__0),
    .in0_0__1(Lift_inst0_out_0__1),
    .in1_0__0(ConcatN_inst2_out_0__0),
    .in1_0__1(ConcatN_inst2_out_0__1),
    .in1_1__0(ConcatN_inst2_out_1__0),
    .in1_1__1(ConcatN_inst2_out_1__1),
    .in1_2__0(ConcatN_inst2_out_2__0),
    .in1_2__1(ConcatN_inst2_out_2__1),
    .out_0__0(ConcatN_inst1_out_0__0),
    .out_0__1(ConcatN_inst1_out_0__1),
    .out_1__0(ConcatN_inst1_out_1__0),
    .out_1__1(ConcatN_inst1_out_1__1),
    .out_2__0(ConcatN_inst1_out_2__0),
    .out_2__1(ConcatN_inst1_out_2__1),
    .out_3__0(ConcatN_inst1_out_3__0),
    .out_3__1(ConcatN_inst1_out_3__1)
);
mantle_concatNArrT__Ns12__t_child_0BitIn_1BitIn2 ConcatN_inst2 (
    .in0_0__0(Lift_inst1_out_0__0),
    .in0_0__1(Lift_inst1_out_0__1),
    .in1_0__0(ConcatN_inst3_out_0__0),
    .in1_0__1(ConcatN_inst3_out_0__1),
    .in1_1__0(ConcatN_inst3_out_1__0),
    .in1_1__1(ConcatN_inst3_out_1__1),
    .out_0__0(ConcatN_inst2_out_0__0),
    .out_0__1(ConcatN_inst2_out_0__1),
    .out_1__0(ConcatN_inst2_out_1__0),
    .out_1__1(ConcatN_inst2_out_1__1),
    .out_2__0(ConcatN_inst2_out_2__0),
    .out_2__1(ConcatN_inst2_out_2__1)
);
mantle_concatNArrT__Ns11__t_child_0BitIn_1BitIn2 ConcatN_inst3 (
    .in0_0__0(Lift_inst2_out_0__0),
    .in0_0__1(Lift_inst2_out_0__1),
    .in1_0__0(ConcatN_inst4_out_0__0),
    .in1_0__1(ConcatN_inst4_out_0__1),
    .out_0__0(ConcatN_inst3_out_0__0),
    .out_0__1(ConcatN_inst3_out_0__1),
    .out_1__0(ConcatN_inst3_out_1__0),
    .out_1__1(ConcatN_inst3_out_1__1)
);
mantle_concatNArrT__Ns1__t_child_0BitIn_1BitIn2 ConcatN_inst4 (
    .in0_0__0(Lift_inst3_out_0__0),
    .in0_0__1(Lift_inst3_out_0__1),
    .out_0__0(ConcatN_inst4_out_0__0),
    .out_0__1(ConcatN_inst4_out_0__1)
);
mantle_concatNArrT__Ns22__t_child_0BitIn_1BitIn2 ConcatN_inst5 (
    .in0_0__0(SlicesBuilder_out0_0__0),
    .in0_0__1(SlicesBuilder_out0_0__1),
    .in0_1__0(SlicesBuilder_out0_1__0),
    .in0_1__1(SlicesBuilder_out0_1__1),
    .in1_0__0(SlicesBuilder_out1_0__0),
    .in1_0__1(SlicesBuilder_out1_0__1),
    .in1_1__0(SlicesBuilder_out1_1__0),
    .in1_1__1(SlicesBuilder_out1_1__1),
    .out_0__0(ConcatN_inst5_out_0__0),
    .out_0__1(ConcatN_inst5_out_0__1),
    .out_1__0(ConcatN_inst5_out_1__0),
    .out_1__1(ConcatN_inst5_out_1__1),
    .out_2__0(ConcatN_inst5_out_2__0),
    .out_2__1(ConcatN_inst5_out_2__1),
    .out_3__0(ConcatN_inst5_out_3__0),
    .out_3__1(ConcatN_inst5_out_3__1)
);
mantle_liftArrT__t_0Bit_1Bit21 Lift_inst0 (
    .in__0(I_1__0),
    .in__1(I_1__1),
    .out_0__0(Lift_inst0_out_0__0),
    .out_0__1(Lift_inst0_out_0__1)
);
mantle_liftArrT__t_0Bit_1Bit21 Lift_inst1 (
    .in__0(I_0__0),
    .in__1(I_0__1),
    .out_0__0(Lift_inst1_out_0__0),
    .out_0__1(Lift_inst1_out_0__1)
);
mantle_liftArrT__t_0Bit_1Bit21 Lift_inst2 (
    .in__0(I_3__0),
    .in__1(I_3__1),
    .out_0__0(Lift_inst2_out_0__0),
    .out_0__1(Lift_inst2_out_0__1)
);
mantle_liftArrT__t_0Bit_1Bit21 Lift_inst3 (
    .in__0(I_2__0),
    .in__1(I_2__1),
    .out_0__0(Lift_inst3_out_0__0),
    .out_0__1(Lift_inst3_out_0__1)
);
mantle_slicesArrT__slices4220__t_0BitIn_1BitIn24 SlicesBuilder (
    .in_0__0(I_0__0),
    .in_0__1(I_0__1),
    .in_1__0(I_1__0),
    .in_1__1(I_1__1),
    .in_2__0(I_2__0),
    .in_2__1(I_2__1),
    .in_3__0(I_3__0),
    .in_3__1(I_3__1),
    .out0_0__0(SlicesBuilder_out0_0__0),
    .out0_0__1(SlicesBuilder_out0_0__1),
    .out0_1__0(SlicesBuilder_out0_1__0),
    .out0_1__1(SlicesBuilder_out0_1__1),
    .out1_0__0(SlicesBuilder_out1_0__0),
    .out1_0__1(SlicesBuilder_out1_0__1),
    .out1_1__0(SlicesBuilder_out1_1__0),
    .out1_1__1(SlicesBuilder_out1_1__1)
);
assign O0_0__0 = I_0__0;
assign O0_0__1 = I_0__1;
assign O0_1__0 = I_1__0;
assign O0_1__1 = I_1__1;
assign O0_2__0 = I_2__0;
assign O0_2__1 = I_2__1;
assign O0_3__0 = I_3__0;
assign O0_3__1 = I_3__1;
assign O1_0__0 = ConcatN_inst0_out_0__0;
assign O1_0__1 = ConcatN_inst0_out_0__1;
assign O1_1__0 = ConcatN_inst0_out_1__0;
assign O1_1__1 = ConcatN_inst0_out_1__1;
assign O1_2__0 = ConcatN_inst0_out_2__0;
assign O1_2__1 = ConcatN_inst0_out_2__1;
assign O1_3__0 = ConcatN_inst0_out_3__0;
assign O1_3__1 = ConcatN_inst0_out_3__1;
assign O2_0__0 = ConcatN_inst1_out_0__0;
assign O2_0__1 = ConcatN_inst1_out_0__1;
assign O2_1__0 = ConcatN_inst1_out_1__0;
assign O2_1__1 = ConcatN_inst1_out_1__1;
assign O2_2__0 = ConcatN_inst1_out_2__0;
assign O2_2__1 = ConcatN_inst1_out_2__1;
assign O2_3__0 = ConcatN_inst1_out_3__0;
assign O2_3__1 = ConcatN_inst1_out_3__1;
assign O3_0__0 = ConcatN_inst5_out_0__0;
assign O3_0__1 = ConcatN_inst5_out_0__1;
assign O3_1__0 = ConcatN_inst5_out_1__0;
assign O3_1__1 = ConcatN_inst5_out_1__1;
assign O3_2__0 = ConcatN_inst5_out_2__0;
assign O3_2__1 = ConcatN_inst5_out_2__1;
assign O3_3__0 = ConcatN_inst5_out_3__0;
assign O3_3__1 = ConcatN_inst5_out_3__1;
endmodule

