module simple_undriven(
  output O
);

  wire _GEN;
  assign O = _GEN;
endmodule

