module simple_custom_verilog_name_custom_name(	// <stdin>:1:1
  input  I,
  output O);

  assign O = I;	// <stdin>:2:5
endmodule

