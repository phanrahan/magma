module LUT(
  input  [1:0]                                         I,
  output struct packed {logic [7:0] x; logic y; }[1:0] O);

  wire [7:0] _tmp = {({{1'h0}, {1'h0}, {1'h0}, {1'h0}})[I], ({{1'h0}, {1'h1}, {1'h1}, {1'h0}})[I], ({{1'h0}, {1'h1}, {1'h0}, {1'h0}})[I], ({{1'h0}, {1'h0}, {1'h0}, {1'h1}})[I], ({{1'h1}, {1'h1}, {1'h1}, {1'h1}})[I], ({{1'h1}, {1'h1}, {1'h0}, {1'h1}})[I], ({{1'h1}, {1'h1}, {1'h1}, {1'h1}})[I], ({{1'h1}, {1'h1}, {1'h1}, {1'h0}})[I]};	// <stdin>:3:14, :4:13, :5:10, :6:10, :7:10, :8:10, :9:10, :10:10, :11:10, :12:10, :13:10, :14:10, :15:11, :16:11, :17:11, :18:11, :19:11, :20:11, :21:11
  wire struct packed {logic [7:0] x; logic y; } _T = '{x: _tmp, y: ({{1'h0}, {1'h1}, {1'h1}, {1'h1}})[I]};	// <stdin>:3:14, :4:13, :5:10, :6:10, :7:10, :8:10, :9:10, :10:10, :11:10, :12:10, :13:10, :14:10, :15:11, :16:11, :17:11, :18:11, :19:11, :20:11, :22:11, :23:11, :24:11
  wire [7:0] _tmp_1 = {({{1'h1}, {1'h1}, {1'h1}, {1'h0}})[I], ({{1'h0}, {1'h1}, {1'h1}, {1'h0}})[I], ({{1'h0}, {1'h0}, {1'h0}, {1'h0}})[I], ({{1'h0}, {1'h0}, {1'h0}, {1'h1}})[I], ({{1'h1}, {1'h0}, {1'h1}, {1'h0}})[I], ({{1'h0}, {1'h0}, {1'h0}, {1'h0}})[I], ({{1'h1}, {1'h1}, {1'h0}, {1'h1}})[I], ({{1'h1}, {1'h1}, {1'h1}, {1'h0}})[I]};	// <stdin>:3:14, :4:13, :25:11, :26:11, :27:11, :28:11, :29:11, :30:11, :31:11, :32:11, :33:11, :34:11, :35:11, :36:11, :37:11, :38:11, :39:11, :40:11, :41:11
  wire struct packed {logic [7:0] x; logic y; } _T_0 = '{x: _tmp_1, y: ({{1'h0}, {1'h0}, {1'h1}, {1'h1}})[I]};	// <stdin>:3:14, :4:13, :25:11, :26:11, :27:11, :28:11, :29:11, :30:11, :31:11, :32:11, :33:11, :34:11, :35:11, :36:11, :37:11, :38:11, :39:11, :40:11, :42:11, :43:11, :44:11
  assign O = {{_T_0}, {_T}};	// <stdin>:45:11, :46:5
endmodule

module complex_lut(
  input  [1:0]                                         a,
  output struct packed {logic [7:0] x; logic y; }[1:0] y);

  LUT LUT_inst0 (	// <stdin>:49:20
    .I (a),
    .O (y)
  );
endmodule

