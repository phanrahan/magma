module test_basic_if_function_call (input [1:0] I, input  S, output  O);
assign O = _O;
endmodule

