module simple_mixed_direction_ports(
  input  [7:0] a_x,
  output [7:0] a_y
);

  assign a_y = a_x;
endmodule

