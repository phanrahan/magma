module coreir_wire #(parameter width = 1) (input [width-1:0] in, output [width-1:0] out);
  assign out = in;
endmodule

module WrappedWire (input I, output O);
wire [0:0] wire_x_O_out;
coreir_wire #(.width(1)) wire_x_O(.in(I), .out(wire_x_O_out));
assign O = wire_x_O_out[0];
endmodule

module Main (input I, output O);
wire wire_x_O_O;
WrappedWire wire_x_O(.I(I), .O(wire_x_O_O));
assign O = wire_x_O_O;
endmodule

