module main (output [0:0] LED, input [0:0] SWITCH);
assign LED = SWITCH;
endmodule

