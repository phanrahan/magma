module basic_if (input [1:0] I, input  S, output  O);
assign O = I[1];
endmodule

