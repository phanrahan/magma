module complex_wire(
  input  [7:0]      I0,
  input             I1,
  input  [3:0][7:0] I2,
  output [7:0]      O0,
  output            O1,
  output [3:0][7:0] O2);

  wire [7:0]  tmp0;	// <stdin>:7:13
  wire        tmp1;	// <stdin>:10:13
  wire [31:0] tmp2;	// <stdin>:78:13

  assign tmp0 = I0;	// <stdin>:8:5
  assign tmp1 = I1;	// <stdin>:11:5
  wire [7:0] _T = I2[2'h0];	// <stdin>:6:14, :13:10
  wire [7:0] _T_0 = I2[2'h0];	// <stdin>:6:14, :15:10
  wire [7:0] _T_1 = I2[2'h0];	// <stdin>:6:14, :17:10
  wire [7:0] _T_2 = I2[2'h0];	// <stdin>:6:14, :19:10
  wire [7:0] _T_3 = I2[2'h0];	// <stdin>:6:14, :21:11
  wire [7:0] _T_4 = I2[2'h0];	// <stdin>:6:14, :23:11
  wire [7:0] _T_5 = I2[2'h0];	// <stdin>:6:14, :25:11
  wire [7:0] _T_6 = I2[2'h0];	// <stdin>:6:14, :27:11
  wire [7:0] _T_7 = I2[2'h1];	// <stdin>:5:14, :29:11
  wire [7:0] _T_8 = I2[2'h1];	// <stdin>:5:14, :31:11
  wire [7:0] _T_9 = I2[2'h1];	// <stdin>:5:14, :33:11
  wire [7:0] _T_10 = I2[2'h1];	// <stdin>:5:14, :35:11
  wire [7:0] _T_11 = I2[2'h1];	// <stdin>:5:14, :37:11
  wire [7:0] _T_12 = I2[2'h1];	// <stdin>:5:14, :39:11
  wire [7:0] _T_13 = I2[2'h1];	// <stdin>:5:14, :41:11
  wire [7:0] _T_14 = I2[2'h1];	// <stdin>:5:14, :43:11
  wire [7:0] _T_15 = I2[2'h2];	// <stdin>:4:15, :45:11
  wire [7:0] _T_16 = I2[2'h2];	// <stdin>:4:15, :47:11
  wire [7:0] _T_17 = I2[2'h2];	// <stdin>:4:15, :49:11
  wire [7:0] _T_18 = I2[2'h2];	// <stdin>:4:15, :51:11
  wire [7:0] _T_19 = I2[2'h2];	// <stdin>:4:15, :53:11
  wire [7:0] _T_20 = I2[2'h2];	// <stdin>:4:15, :55:11
  wire [7:0] _T_21 = I2[2'h2];	// <stdin>:4:15, :57:11
  wire [7:0] _T_22 = I2[2'h2];	// <stdin>:4:15, :59:11
  wire [7:0] _T_23 = I2[2'h3];	// <stdin>:3:15, :61:11
  wire [7:0] _T_24 = I2[2'h3];	// <stdin>:3:15, :63:11
  wire [7:0] _T_25 = I2[2'h3];	// <stdin>:3:15, :65:11
  wire [7:0] _T_26 = I2[2'h3];	// <stdin>:3:15, :67:11
  wire [7:0] _T_27 = I2[2'h3];	// <stdin>:3:15, :69:11
  wire [7:0] _T_28 = I2[2'h3];	// <stdin>:3:15, :71:11
  wire [7:0] _T_29 = I2[2'h3];	// <stdin>:3:15, :73:11
  wire [7:0] _T_30 = I2[2'h3];	// <stdin>:3:15, :75:11
  assign tmp2 = {_T_30[7], _T_29[6], _T_28[5], _T_27[4], _T_26[3], _T_25[2], _T_24[1], _T_23[0], _T_22[7], _T_21[6], _T_20[5], _T_19[4], _T_18[3], _T_17[2], _T_16[1], _T_15[0], _T_14[7], _T_13[6], _T_12[5], _T_11[4], _T_10[3], _T_9[2], _T_8[1], _T_7[0], _T_6[7], _T_5[6], _T_4[5], _T_3[4], _T_2[3], _T_1[2], _T_0[1], _T[0]};	// <stdin>:14:10, :16:10, :18:10, :20:10, :22:11, :24:11, :26:11, :28:11, :30:11, :32:11, :34:11, :36:11, :38:11, :40:11, :42:11, :44:11, :46:11, :48:11, :50:11, :52:11, :54:11, :56:11, :58:11, :60:11, :62:11, :64:11, :66:11, :68:11, :70:11, :72:11, :74:11, :76:11, :77:11, :79:5
  wire [31:0] _T_31 = tmp2;	// <stdin>:80:11
  assign O0 = tmp0;	// <stdin>:9:10, :86:5
  assign O1 = tmp1;	// <stdin>:12:10, :86:5
  assign O2 = {{_T_31[31:24]}, {_T_31[23:16]}, {_T_31[15:8]}, {_T_31[7:0]}};	// <stdin>:81:11, :82:11, :83:11, :84:11, :85:11, :86:5
endmodule

