module mod3 #(parameter KRATOS_INSTANCE_ID = 16'b1)
(
    input I
);

endmodule   // mod
