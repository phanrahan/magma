module Bar (
    input I,
    output O
);
assign O = I;
endmodule

