module if_statement_nested (input [3:0] I, input [1:0] S, output  O);
assign O = I[3];
endmodule

