module feedthrough(
  input  I,
  output O
);

  assign O = I;
endmodule

