module simple_length_one_bits(	// <stdin>:1:1
  input  I,
  output O);

  assign O = I;	// <stdin>:3:5
endmodule

