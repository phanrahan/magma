module main (output [1:0] O);
assign O = 2'd2';
endmodule

