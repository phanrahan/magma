module simple_magma_protocol(
  input  [7:0] I,
  output [7:0] O
);

  assign O = I;
endmodule

