module simple_undriven(	// <stdin>:1:1
  output O);

  wire _T;	// <stdin>:2:10

  assign O = _T;	// <stdin>:3:10, :4:5
endmodule

