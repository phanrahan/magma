module bar_foo_OtherCircuit (
    output [19:0] x_y [0:0]
);
endmodule
