module mod4 #(parameter KRATOS_INSTANCE_ID = 13'o742)
(
    input I
);

endmodule   // mod
