module if_statement_nested (input [3:0] I_0, input [1:0] S_0, output  O);
assign O = I_0[3];
endmodule

