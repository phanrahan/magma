module simple_inline_verilog(
  input  I,
  output O);

  
  	// This is 'a' "comment".	// <stdin>:4:5
  assign O = I;	// <stdin>:5:5
endmodule

