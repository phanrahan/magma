module Main (input I, output O);
assign O = I;
endmodule

