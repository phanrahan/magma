module mod3 #(parameter KRATOS_INSTANCE_ID = 16'b10111)
(
    input I
);

endmodule   // mod
