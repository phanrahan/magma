module BasicALU(	// <stdin>:1:1
  input  [3:0] a, b, opcode,
  output [3:0] out);

  wire [1:0][3:0] _T = {{{3'h0, a == b}}, {{3'h0, a < b}}};	// <stdin>:2:10, :6:10, :7:10, :11:10, :14:11
  wire [1:0][3:0] _T_0 = {{_T[opcode == 4'h8]}, {a - b}};	// <stdin>:12:11, :13:11, :15:11, :16:11, :19:11
  wire [1:0][3:0] _T_1 = {{_T_0[opcode == 4'h7]}, {a + b}};	// <stdin>:17:11, :18:11, :20:11, :21:11, :24:11
  wire [1:0][3:0] _T_2 = {{_T_1[opcode == 4'h6]}, {a - 4'h4}};	// <stdin>:22:11, :23:11, :25:11, :27:11, :30:11
  wire [1:0][3:0] _T_3 = {{_T_2[opcode == 4'h5]}, {a + 4'h4}};	// <stdin>:28:11, :29:11, :31:11, :32:11, :33:11, :36:11
  wire [1:0][3:0] _T_4 = {{_T_3[opcode == 4'h4]}, {a - 4'h1}};	// <stdin>:32:11, :35:11, :37:11, :39:11, :42:11
  wire [1:0][3:0] _T_5 = {{_T_4[opcode == 4'h3]}, {a + 4'h1}};	// <stdin>:40:11, :41:11, :43:11, :44:11, :45:11, :48:11
  wire [1:0][3:0] _T_6 = {{_T_5[opcode == 4'h2]}, {b}};	// <stdin>:46:11, :47:11, :49:11, :52:11
  wire [1:0][3:0] _T_7 = {{_T_6[opcode == 4'h1]}, {a}};	// <stdin>:44:11, :51:11, :53:11, :56:11
  assign out = _T_7[opcode == 4'h0];	// <stdin>:54:11, :55:11, :57:11, :58:5
endmodule

