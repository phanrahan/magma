module return_magma_named_tuple (input [1:0] I_0, output  O_x, output  O_y);
assign O_x = I_0[0];
assign O_y = I_0[1];
endmodule

