module complex_aggregates_nested_array(	// <stdin>:1:1
  input  [1:0][2:0][3:0] a,
  output [1:0][2:0][3:0] y);

  wire [2:0][3:0] _T = a[1'h0];	// <stdin>:2:10, :3:10
  wire [3:0] _T_0 = _T[2'h0];	// <stdin>:4:10, :5:10
  wire _T_1 = _T_0[0];	// <stdin>:6:10
  wire [2:0][3:0] _T_2 = a[1'h1];	// <stdin>:7:10, :8:10
  wire [3:0] _T_3 = _T_2[2'h2];	// <stdin>:9:10, :10:10
  wire _T_4 = _T_3[3];	// <stdin>:11:10
  wire _T_5 = _T_0[1];	// <stdin>:13:11
  wire _T_6 = _T_3[2];	// <stdin>:14:11
  wire _T_7 = _T_0[2];	// <stdin>:16:11
  wire _T_8 = _T_3[1];	// <stdin>:17:11
  wire _T_9 = _T_0[3];	// <stdin>:19:11
  wire _T_10 = _T_3[0];	// <stdin>:20:11
  wire [3:0] _T_11 = _T[2'h1];	// <stdin>:23:11, :24:11
  wire _T_12 = _T_11[0];	// <stdin>:25:11
  wire [3:0] _T_13 = _T_2[2'h1];	// <stdin>:23:11, :26:11
  wire _T_14 = _T_13[3];	// <stdin>:27:11
  wire _T_15 = _T_11[1];	// <stdin>:29:11
  wire _T_16 = _T_13[2];	// <stdin>:30:11
  wire _T_17 = _T_11[2];	// <stdin>:32:11
  wire _T_18 = _T_13[1];	// <stdin>:33:11
  wire _T_19 = _T_11[3];	// <stdin>:35:11
  wire _T_20 = _T_13[0];	// <stdin>:36:11
  wire [3:0] _T_21 = _T[2'h2];	// <stdin>:9:10, :39:11
  wire _T_22 = _T_21[0];	// <stdin>:40:11
  wire [3:0] _T_23 = _T_2[2'h0];	// <stdin>:4:10, :41:11
  wire _T_24 = _T_23[3];	// <stdin>:42:11
  wire _T_25 = _T_21[1];	// <stdin>:44:11
  wire _T_26 = _T_23[2];	// <stdin>:45:11
  wire _T_27 = _T_21[2];	// <stdin>:47:11
  wire _T_28 = _T_23[1];	// <stdin>:48:11
  wire _T_29 = _T_21[3];	// <stdin>:50:11
  wire _T_30 = _T_23[0];	// <stdin>:51:11
  assign y = {{{{{_T_4 | _T_1, _T_6 | _T_5, _T_8 | _T_7, _T_10 | _T_9}}, {{_T_14 | _T_12, _T_16 | _T_15,
                _T_18 | _T_17, _T_20 | _T_19}}, {{_T_24 | _T_22, _T_26 | _T_25, _T_28 | _T_27, _T_30 |
                _T_29}}}}, {{{{_T_29 | _T_30, _T_27 | _T_28, _T_25 | _T_26, _T_22 | _T_24}}, {{_T_19 |
                _T_20, _T_17 | _T_18, _T_15 | _T_16, _T_12 | _T_14}}, {{_T_9 | _T_10, _T_7 | _T_8, _T_5 |
                _T_6, _T_1 | _T_4}}}}};	// <stdin>:12:11, :15:11, :18:11, :21:11, :22:11, :28:11, :31:11, :34:11, :37:11, :38:11, :43:11, :46:11, :49:11, :52:11, :53:11, :54:11, :55:11, :56:11, :57:11, :58:11, :59:11, :60:11, :61:11, :62:11, :63:11, :64:11, :65:11, :66:11, :67:11, :68:11, :69:11, :70:11, :71:11, :72:5
endmodule

