module test_reduce_and_ (
    input [4:0] I,
    output O
);
assign O = & I;
endmodule

