module simple_clock_cast(
  input  I,
  output O
);

  assign O = I;
endmodule

