module main (output [1:0] O);
assign O = {1'b1,1'b0};
endmodule

