module mantle_wire__type_0Bit_1Bit23 (
    input in_0__0,
    input [1:0] in_0__1,
    input in_1__0,
    input [1:0] in_1__1,
    input in_2__0,
    input [1:0] in_2__1,
    output out_0__0,
    output [1:0] out_0__1,
    output out_1__0,
    output [1:0] out_1__1,
    output out_2__0,
    output [1:0] out_2__1
);
assign out_0__0 = in_0__0;
assign out_0__1 = in_0__1;
assign out_1__0 = in_1__0;
assign out_1__1 = in_1__1;
assign out_2__0 = in_2__0;
assign out_2__1 = in_2__1;
endmodule

module mantle_wire__type_0Bit_1Bit22 (
    input in_0__0,
    input [1:0] in_0__1,
    input in_1__0,
    input [1:0] in_1__1,
    output out_0__0,
    output [1:0] out_0__1,
    output out_1__0,
    output [1:0] out_1__1
);
assign out_0__0 = in_0__0;
assign out_0__1 = in_0__1;
assign out_1__0 = in_1__0;
assign out_1__1 = in_1__1;
endmodule

module mantle_wire__type_0Bit_1Bit21 (
    input in_0__0,
    input [1:0] in_0__1,
    output out_0__0,
    output [1:0] out_0__1
);
assign out_0__0 = in_0__0;
assign out_0__1 = in_0__1;
endmodule

module mantle_wire__type_0Bit_1Bit2 (
    input in__0,
    input [1:0] in__1,
    output out__0,
    output [1:0] out__1
);
assign out__0 = in__0;
assign out__1 = in__1;
endmodule

module mantle_liftArrT__t_0Bit_1Bit21 (
    input in__0,
    input [1:0] in__1,
    output out_0__0,
    output [1:0] out_0__1
);
assign out_0__0 = in__0;
assign out_0__1 = in__1;
endmodule

module mantle_getArrT__i3__t_0BitIn_1BitIn24 (
    input in_0__0,
    input [1:0] in_0__1,
    input in_1__0,
    input [1:0] in_1__1,
    input in_2__0,
    input [1:0] in_2__1,
    input in_3__0,
    input [1:0] in_3__1,
    output out__0,
    output [1:0] out__1
);
assign out__0 = in_3__0;
assign out__1 = in_3__1;
endmodule

module mantle_getArrT__i2__t_0BitIn_1BitIn24 (
    input in_0__0,
    input [1:0] in_0__1,
    input in_1__0,
    input [1:0] in_1__1,
    input in_2__0,
    input [1:0] in_2__1,
    input in_3__0,
    input [1:0] in_3__1,
    output out__0,
    output [1:0] out__1
);
assign out__0 = in_2__0;
assign out__1 = in_2__1;
endmodule

module mantle_getArrT__i1__t_0BitIn_1BitIn24 (
    input in_0__0,
    input [1:0] in_0__1,
    input in_1__0,
    input [1:0] in_1__1,
    input in_2__0,
    input [1:0] in_2__1,
    input in_3__0,
    input [1:0] in_3__1,
    output out__0,
    output [1:0] out__1
);
assign out__0 = in_1__0;
assign out__1 = in_1__1;
endmodule

module mantle_getArrT__i0__t_0BitIn_1BitIn24 (
    input in_0__0,
    input [1:0] in_0__1,
    input in_1__0,
    input [1:0] in_1__1,
    input in_2__0,
    input [1:0] in_2__1,
    input in_3__0,
    input [1:0] in_3__1,
    output out__0,
    output [1:0] out__1
);
assign out__0 = in_0__0;
assign out__1 = in_0__1;
endmodule

module mantle_concatArrT__t0_0BitIn_1BitIn21__t1_0BitIn_1BitIn23 (
    input in0_0__0,
    input [1:0] in0_0__1,
    input in1_0__0,
    input [1:0] in1_0__1,
    input in1_1__0,
    input [1:0] in1_1__1,
    input in1_2__0,
    input [1:0] in1_2__1,
    output out_0__0,
    output [1:0] out_0__1,
    output out_1__0,
    output [1:0] out_1__1,
    output out_2__0,
    output [1:0] out_2__1,
    output out_3__0,
    output [1:0] out_3__1
);
assign out_0__0 = in0_0__0;
assign out_0__1 = in0_0__1;
assign out_1__0 = in1_0__0;
assign out_1__1 = in1_0__1;
assign out_2__0 = in1_1__0;
assign out_2__1 = in1_1__1;
assign out_3__0 = in1_2__0;
assign out_3__1 = in1_2__1;
endmodule

module mantle_concatArrT__t0_0BitIn_1BitIn21__t1_0BitIn_1BitIn22 (
    input in0_0__0,
    input [1:0] in0_0__1,
    input in1_0__0,
    input [1:0] in1_0__1,
    input in1_1__0,
    input [1:0] in1_1__1,
    output out_0__0,
    output [1:0] out_0__1,
    output out_1__0,
    output [1:0] out_1__1,
    output out_2__0,
    output [1:0] out_2__1
);
assign out_0__0 = in0_0__0;
assign out_0__1 = in0_0__1;
assign out_1__0 = in1_0__0;
assign out_1__1 = in1_0__1;
assign out_2__0 = in1_1__0;
assign out_2__1 = in1_1__1;
endmodule

module mantle_concatArrT__t0_0BitIn_1BitIn21__t1_0BitIn_1BitIn21 (
    input in0_0__0,
    input [1:0] in0_0__1,
    input in1_0__0,
    input [1:0] in1_0__1,
    output out_0__0,
    output [1:0] out_0__1,
    output out_1__0,
    output [1:0] out_1__1
);
assign out_0__0 = in0_0__0;
assign out_0__1 = in0_0__1;
assign out_1__0 = in1_0__0;
assign out_1__1 = in1_0__1;
endmodule

module Foo (
    input I_0__0,
    input [1:0] I_0__1,
    input I_1__0,
    input [1:0] I_1__1,
    input I_2__0,
    input [1:0] I_2__1,
    input I_3__0,
    input [1:0] I_3__1,
    output O_0__0,
    output [1:0] O_0__1,
    output O_1__0,
    output [1:0] O_1__1,
    output O_2__0,
    output [1:0] O_2__1,
    output O_3__0,
    output [1:0] O_3__1
);
wire Concat_inst0_out_0__0;
wire [1:0] Concat_inst0_out_0__1;
wire Concat_inst0_out_1__0;
wire [1:0] Concat_inst0_out_1__1;
wire Concat_inst0_out_2__0;
wire [1:0] Concat_inst0_out_2__1;
wire Concat_inst0_out_3__0;
wire [1:0] Concat_inst0_out_3__1;
wire Concat_inst1_out_0__0;
wire [1:0] Concat_inst1_out_0__1;
wire Concat_inst1_out_1__0;
wire [1:0] Concat_inst1_out_1__1;
wire Concat_inst1_out_2__0;
wire [1:0] Concat_inst1_out_2__1;
wire Concat_inst2_out_0__0;
wire [1:0] Concat_inst2_out_0__1;
wire Concat_inst2_out_1__0;
wire [1:0] Concat_inst2_out_1__1;
wire Index_inst0_out__0;
wire [1:0] Index_inst0_out__1;
wire Index_inst1_out__0;
wire [1:0] Index_inst1_out__1;
wire Index_inst2_out__0;
wire [1:0] Index_inst2_out__1;
wire Index_inst3_out__0;
wire [1:0] Index_inst3_out__1;
wire Index_inst4_out__0;
wire [1:0] Index_inst4_out__1;
wire Index_inst5_out__0;
wire [1:0] Index_inst5_out__1;
wire Index_inst6_out__0;
wire [1:0] Index_inst6_out__1;
wire Index_inst7_out__0;
wire [1:0] Index_inst7_out__1;
wire Lift_inst0_out_0__0;
wire [1:0] Lift_inst0_out_0__1;
wire Lift_inst1_out_0__0;
wire [1:0] Lift_inst1_out_0__1;
wire Lift_inst2_out_0__0;
wire [1:0] Lift_inst2_out_0__1;
wire Lift_inst3_out_0__0;
wire [1:0] Lift_inst3_out_0__1;
wire Wire_inst0_out__0;
wire [1:0] Wire_inst0_out__1;
wire Wire_inst1_out_0__0;
wire [1:0] Wire_inst1_out_0__1;
wire Wire_inst1_out_1__0;
wire [1:0] Wire_inst1_out_1__1;
wire Wire_inst1_out_2__0;
wire [1:0] Wire_inst1_out_2__1;
wire Wire_inst2_out__0;
wire [1:0] Wire_inst2_out__1;
wire Wire_inst3_out_0__0;
wire [1:0] Wire_inst3_out_0__1;
wire Wire_inst3_out_1__0;
wire [1:0] Wire_inst3_out_1__1;
wire Wire_inst4_out__0;
wire [1:0] Wire_inst4_out__1;
wire Wire_inst5_out_0__0;
wire [1:0] Wire_inst5_out_0__1;
wire Wire_inst6_out__0;
wire [1:0] Wire_inst6_out__1;
mantle_concatArrT__t0_0BitIn_1BitIn21__t1_0BitIn_1BitIn23 Concat_inst0 (
    .in0_0__0(Lift_inst0_out_0__0),
    .in0_0__1(Lift_inst0_out_0__1),
    .in1_0__0(Wire_inst1_out_0__0),
    .in1_0__1(Wire_inst1_out_0__1),
    .in1_1__0(Wire_inst1_out_1__0),
    .in1_1__1(Wire_inst1_out_1__1),
    .in1_2__0(Wire_inst1_out_2__0),
    .in1_2__1(Wire_inst1_out_2__1),
    .out_0__0(Concat_inst0_out_0__0),
    .out_0__1(Concat_inst0_out_0__1),
    .out_1__0(Concat_inst0_out_1__0),
    .out_1__1(Concat_inst0_out_1__1),
    .out_2__0(Concat_inst0_out_2__0),
    .out_2__1(Concat_inst0_out_2__1),
    .out_3__0(Concat_inst0_out_3__0),
    .out_3__1(Concat_inst0_out_3__1)
);
mantle_concatArrT__t0_0BitIn_1BitIn21__t1_0BitIn_1BitIn22 Concat_inst1 (
    .in0_0__0(Lift_inst1_out_0__0),
    .in0_0__1(Lift_inst1_out_0__1),
    .in1_0__0(Wire_inst3_out_0__0),
    .in1_0__1(Wire_inst3_out_0__1),
    .in1_1__0(Wire_inst3_out_1__0),
    .in1_1__1(Wire_inst3_out_1__1),
    .out_0__0(Concat_inst1_out_0__0),
    .out_0__1(Concat_inst1_out_0__1),
    .out_1__0(Concat_inst1_out_1__0),
    .out_1__1(Concat_inst1_out_1__1),
    .out_2__0(Concat_inst1_out_2__0),
    .out_2__1(Concat_inst1_out_2__1)
);
mantle_concatArrT__t0_0BitIn_1BitIn21__t1_0BitIn_1BitIn21 Concat_inst2 (
    .in0_0__0(Lift_inst2_out_0__0),
    .in0_0__1(Lift_inst2_out_0__1),
    .in1_0__0(Wire_inst5_out_0__0),
    .in1_0__1(Wire_inst5_out_0__1),
    .out_0__0(Concat_inst2_out_0__0),
    .out_0__1(Concat_inst2_out_0__1),
    .out_1__0(Concat_inst2_out_1__0),
    .out_1__1(Concat_inst2_out_1__1)
);
mantle_getArrT__i3__t_0BitIn_1BitIn24 Index_inst0 (
    .in_0__0(I_0__0),
    .in_0__1(I_0__1),
    .in_1__0(I_1__0),
    .in_1__1(I_1__1),
    .in_2__0(I_2__0),
    .in_2__1(I_2__1),
    .in_3__0(I_3__0),
    .in_3__1(I_3__1),
    .out__0(Index_inst0_out__0),
    .out__1(Index_inst0_out__1)
);
mantle_getArrT__i0__t_0BitIn_1BitIn24 Index_inst1 (
    .in_0__0(I_0__0),
    .in_0__1(I_0__1),
    .in_1__0(I_1__0),
    .in_1__1(I_1__1),
    .in_2__0(I_2__0),
    .in_2__1(I_2__1),
    .in_3__0(I_3__0),
    .in_3__1(I_3__1),
    .out__0(Index_inst1_out__0),
    .out__1(Index_inst1_out__1)
);
mantle_getArrT__i2__t_0BitIn_1BitIn24 Index_inst2 (
    .in_0__0(I_0__0),
    .in_0__1(I_0__1),
    .in_1__0(I_1__0),
    .in_1__1(I_1__1),
    .in_2__0(I_2__0),
    .in_2__1(I_2__1),
    .in_3__0(I_3__0),
    .in_3__1(I_3__1),
    .out__0(Index_inst2_out__0),
    .out__1(Index_inst2_out__1)
);
mantle_getArrT__i1__t_0BitIn_1BitIn24 Index_inst3 (
    .in_0__0(I_0__0),
    .in_0__1(I_0__1),
    .in_1__0(I_1__0),
    .in_1__1(I_1__1),
    .in_2__0(I_2__0),
    .in_2__1(I_2__1),
    .in_3__0(I_3__0),
    .in_3__1(I_3__1),
    .out__0(Index_inst3_out__0),
    .out__1(Index_inst3_out__1)
);
mantle_getArrT__i1__t_0BitIn_1BitIn24 Index_inst4 (
    .in_0__0(I_0__0),
    .in_0__1(I_0__1),
    .in_1__0(I_1__0),
    .in_1__1(I_1__1),
    .in_2__0(I_2__0),
    .in_2__1(I_2__1),
    .in_3__0(I_3__0),
    .in_3__1(I_3__1),
    .out__0(Index_inst4_out__0),
    .out__1(Index_inst4_out__1)
);
mantle_getArrT__i2__t_0BitIn_1BitIn24 Index_inst5 (
    .in_0__0(I_0__0),
    .in_0__1(I_0__1),
    .in_1__0(I_1__0),
    .in_1__1(I_1__1),
    .in_2__0(I_2__0),
    .in_2__1(I_2__1),
    .in_3__0(I_3__0),
    .in_3__1(I_3__1),
    .out__0(Index_inst5_out__0),
    .out__1(Index_inst5_out__1)
);
mantle_getArrT__i0__t_0BitIn_1BitIn24 Index_inst6 (
    .in_0__0(I_0__0),
    .in_0__1(I_0__1),
    .in_1__0(I_1__0),
    .in_1__1(I_1__1),
    .in_2__0(I_2__0),
    .in_2__1(I_2__1),
    .in_3__0(I_3__0),
    .in_3__1(I_3__1),
    .out__0(Index_inst6_out__0),
    .out__1(Index_inst6_out__1)
);
mantle_getArrT__i3__t_0BitIn_1BitIn24 Index_inst7 (
    .in_0__0(I_0__0),
    .in_0__1(I_0__1),
    .in_1__0(I_1__0),
    .in_1__1(I_1__1),
    .in_2__0(I_2__0),
    .in_2__1(I_2__1),
    .in_3__0(I_3__0),
    .in_3__1(I_3__1),
    .out__0(Index_inst7_out__0),
    .out__1(Index_inst7_out__1)
);
mantle_liftArrT__t_0Bit_1Bit21 Lift_inst0 (
    .in__0(Wire_inst0_out__0),
    .in__1(Wire_inst0_out__1),
    .out_0__0(Lift_inst0_out_0__0),
    .out_0__1(Lift_inst0_out_0__1)
);
mantle_liftArrT__t_0Bit_1Bit21 Lift_inst1 (
    .in__0(Wire_inst2_out__0),
    .in__1(Wire_inst2_out__1),
    .out_0__0(Lift_inst1_out_0__0),
    .out_0__1(Lift_inst1_out_0__1)
);
mantle_liftArrT__t_0Bit_1Bit21 Lift_inst2 (
    .in__0(Wire_inst4_out__0),
    .in__1(Wire_inst4_out__1),
    .out_0__0(Lift_inst2_out_0__0),
    .out_0__1(Lift_inst2_out_0__1)
);
mantle_liftArrT__t_0Bit_1Bit21 Lift_inst3 (
    .in__0(Wire_inst6_out__0),
    .in__1(Wire_inst6_out__1),
    .out_0__0(Lift_inst3_out_0__0),
    .out_0__1(Lift_inst3_out_0__1)
);
mantle_wire__type_0Bit_1Bit2 Wire_inst0 (
    .in__0(Index_inst0_out__0),
    .in__1(Index_inst1_out__1),
    .out__0(Wire_inst0_out__0),
    .out__1(Wire_inst0_out__1)
);
mantle_wire__type_0Bit_1Bit23 Wire_inst1 (
    .in_0__0(Concat_inst1_out_0__0),
    .in_0__1(Concat_inst1_out_0__1),
    .in_1__0(Concat_inst1_out_1__0),
    .in_1__1(Concat_inst1_out_1__1),
    .in_2__0(Concat_inst1_out_2__0),
    .in_2__1(Concat_inst1_out_2__1),
    .out_0__0(Wire_inst1_out_0__0),
    .out_0__1(Wire_inst1_out_0__1),
    .out_1__0(Wire_inst1_out_1__0),
    .out_1__1(Wire_inst1_out_1__1),
    .out_2__0(Wire_inst1_out_2__0),
    .out_2__1(Wire_inst1_out_2__1)
);
mantle_wire__type_0Bit_1Bit2 Wire_inst2 (
    .in__0(Index_inst2_out__0),
    .in__1(Index_inst3_out__1),
    .out__0(Wire_inst2_out__0),
    .out__1(Wire_inst2_out__1)
);
mantle_wire__type_0Bit_1Bit22 Wire_inst3 (
    .in_0__0(Concat_inst2_out_0__0),
    .in_0__1(Concat_inst2_out_0__1),
    .in_1__0(Concat_inst2_out_1__0),
    .in_1__1(Concat_inst2_out_1__1),
    .out_0__0(Wire_inst3_out_0__0),
    .out_0__1(Wire_inst3_out_0__1),
    .out_1__0(Wire_inst3_out_1__0),
    .out_1__1(Wire_inst3_out_1__1)
);
mantle_wire__type_0Bit_1Bit2 Wire_inst4 (
    .in__0(Index_inst4_out__0),
    .in__1(Index_inst5_out__1),
    .out__0(Wire_inst4_out__0),
    .out__1(Wire_inst4_out__1)
);
mantle_wire__type_0Bit_1Bit21 Wire_inst5 (
    .in_0__0(Lift_inst3_out_0__0),
    .in_0__1(Lift_inst3_out_0__1),
    .out_0__0(Wire_inst5_out_0__0),
    .out_0__1(Wire_inst5_out_0__1)
);
mantle_wire__type_0Bit_1Bit2 Wire_inst6 (
    .in__0(Index_inst6_out__0),
    .in__1(Index_inst7_out__1),
    .out__0(Wire_inst6_out__0),
    .out__1(Wire_inst6_out__1)
);
assign O_0__0 = Concat_inst0_out_0__0;
assign O_0__1 = Concat_inst0_out_0__1;
assign O_1__0 = Concat_inst0_out_1__0;
assign O_1__1 = Concat_inst0_out_1__1;
assign O_2__0 = Concat_inst0_out_2__0;
assign O_2__1 = Concat_inst0_out_2__1;
assign O_3__0 = Concat_inst0_out_3__0;
assign O_3__1 = Concat_inst0_out_3__1;
endmodule

