module mod2 #(parameter KRATOS_INSTANCE_ID = 24'sd2)
(
    input I
);

endmodule   // mod
