module main (output  O);
assign O = 1'b1;
endmodule

